// Core3.v

// Generated using ACDS version 13.0sp1 232 at 2021.05.28.02:37:29

`timescale 1 ps / 1 ps
module Core3 (
		input  wire        clk_clk,                               //                            clk.clk
		output wire [17:0] red_leds_external_connection_export,   //   red_leds_external_connection.export
		output wire [7:0]  green_leds_external_connection_export, // green_leds_external_connection.export
		input  wire [17:0] switches_external_connection_export,   //   switches_external_connection.export
		input  wire        reset_reset_n                          //                          reset.reset_n
	);

	wire         cpu_0_instruction_master_waitrequest;                                                                     // cpu_0_instruction_master_translator:av_waitrequest -> cpu_0:i_waitrequest
	wire  [17:0] cpu_0_instruction_master_address;                                                                         // cpu_0:i_address -> cpu_0_instruction_master_translator:av_address
	wire         cpu_0_instruction_master_read;                                                                            // cpu_0:i_read -> cpu_0_instruction_master_translator:av_read
	wire  [31:0] cpu_0_instruction_master_readdata;                                                                        // cpu_0_instruction_master_translator:av_readdata -> cpu_0:i_readdata
	wire         cpu_0_data_master_waitrequest;                                                                            // cpu_0_data_master_translator:av_waitrequest -> cpu_0:d_waitrequest
	wire  [31:0] cpu_0_data_master_writedata;                                                                              // cpu_0:d_writedata -> cpu_0_data_master_translator:av_writedata
	wire  [17:0] cpu_0_data_master_address;                                                                                // cpu_0:d_address -> cpu_0_data_master_translator:av_address
	wire         cpu_0_data_master_write;                                                                                  // cpu_0:d_write -> cpu_0_data_master_translator:av_write
	wire         cpu_0_data_master_read;                                                                                   // cpu_0:d_read -> cpu_0_data_master_translator:av_read
	wire  [31:0] cpu_0_data_master_readdata;                                                                               // cpu_0_data_master_translator:av_readdata -> cpu_0:d_readdata
	wire         cpu_0_data_master_debugaccess;                                                                            // cpu_0:jtag_debug_module_debugaccess_to_roms -> cpu_0_data_master_translator:av_debugaccess
	wire   [3:0] cpu_0_data_master_byteenable;                                                                             // cpu_0:d_byteenable -> cpu_0_data_master_translator:av_byteenable
	wire         cpu_1_data_master_waitrequest;                                                                            // cpu_1_data_master_translator:av_waitrequest -> cpu_1:d_waitrequest
	wire  [31:0] cpu_1_data_master_writedata;                                                                              // cpu_1:d_writedata -> cpu_1_data_master_translator:av_writedata
	wire  [17:0] cpu_1_data_master_address;                                                                                // cpu_1:d_address -> cpu_1_data_master_translator:av_address
	wire         cpu_1_data_master_write;                                                                                  // cpu_1:d_write -> cpu_1_data_master_translator:av_write
	wire         cpu_1_data_master_read;                                                                                   // cpu_1:d_read -> cpu_1_data_master_translator:av_read
	wire  [31:0] cpu_1_data_master_readdata;                                                                               // cpu_1_data_master_translator:av_readdata -> cpu_1:d_readdata
	wire         cpu_1_data_master_debugaccess;                                                                            // cpu_1:jtag_debug_module_debugaccess_to_roms -> cpu_1_data_master_translator:av_debugaccess
	wire   [3:0] cpu_1_data_master_byteenable;                                                                             // cpu_1:d_byteenable -> cpu_1_data_master_translator:av_byteenable
	wire         cpu_2_data_master_waitrequest;                                                                            // cpu_2_data_master_translator:av_waitrequest -> cpu_2:d_waitrequest
	wire  [31:0] cpu_2_data_master_writedata;                                                                              // cpu_2:d_writedata -> cpu_2_data_master_translator:av_writedata
	wire  [17:0] cpu_2_data_master_address;                                                                                // cpu_2:d_address -> cpu_2_data_master_translator:av_address
	wire         cpu_2_data_master_write;                                                                                  // cpu_2:d_write -> cpu_2_data_master_translator:av_write
	wire         cpu_2_data_master_read;                                                                                   // cpu_2:d_read -> cpu_2_data_master_translator:av_read
	wire  [31:0] cpu_2_data_master_readdata;                                                                               // cpu_2_data_master_translator:av_readdata -> cpu_2:d_readdata
	wire         cpu_2_data_master_debugaccess;                                                                            // cpu_2:jtag_debug_module_debugaccess_to_roms -> cpu_2_data_master_translator:av_debugaccess
	wire   [3:0] cpu_2_data_master_byteenable;                                                                             // cpu_2:d_byteenable -> cpu_2_data_master_translator:av_byteenable
	wire         cpu_1_instruction_master_waitrequest;                                                                     // cpu_1_instruction_master_translator:av_waitrequest -> cpu_1:i_waitrequest
	wire  [17:0] cpu_1_instruction_master_address;                                                                         // cpu_1:i_address -> cpu_1_instruction_master_translator:av_address
	wire         cpu_1_instruction_master_read;                                                                            // cpu_1:i_read -> cpu_1_instruction_master_translator:av_read
	wire  [31:0] cpu_1_instruction_master_readdata;                                                                        // cpu_1_instruction_master_translator:av_readdata -> cpu_1:i_readdata
	wire         cpu_2_instruction_master_waitrequest;                                                                     // cpu_2_instruction_master_translator:av_waitrequest -> cpu_2:i_waitrequest
	wire  [17:0] cpu_2_instruction_master_address;                                                                         // cpu_2:i_address -> cpu_2_instruction_master_translator:av_address
	wire         cpu_2_instruction_master_read;                                                                            // cpu_2:i_read -> cpu_2_instruction_master_translator:av_read
	wire  [31:0] cpu_2_instruction_master_readdata;                                                                        // cpu_2_instruction_master_translator:av_readdata -> cpu_2:i_readdata
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                       // cpu_0:jtag_debug_module_waitrequest -> cpu_0_jtag_debug_module_translator:av_waitrequest
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                         // cpu_0_jtag_debug_module_translator:av_writedata -> cpu_0:jtag_debug_module_writedata
	wire   [8:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                                           // cpu_0_jtag_debug_module_translator:av_address -> cpu_0:jtag_debug_module_address
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                             // cpu_0_jtag_debug_module_translator:av_write -> cpu_0:jtag_debug_module_write
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_read;                                              // cpu_0_jtag_debug_module_translator:av_read -> cpu_0:jtag_debug_module_read
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                          // cpu_0:jtag_debug_module_readdata -> cpu_0_jtag_debug_module_translator:av_readdata
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                       // cpu_0_jtag_debug_module_translator:av_debugaccess -> cpu_0:jtag_debug_module_debugaccess
	wire   [3:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                        // cpu_0_jtag_debug_module_translator:av_byteenable -> cpu_0:jtag_debug_module_byteenable
	wire  [31:0] onchip_memory_0_s1_translator_avalon_anti_slave_0_writedata;                                              // onchip_memory_0_s1_translator:av_writedata -> onchip_memory_0:writedata
	wire  [12:0] onchip_memory_0_s1_translator_avalon_anti_slave_0_address;                                                // onchip_memory_0_s1_translator:av_address -> onchip_memory_0:address
	wire         onchip_memory_0_s1_translator_avalon_anti_slave_0_chipselect;                                             // onchip_memory_0_s1_translator:av_chipselect -> onchip_memory_0:chipselect
	wire         onchip_memory_0_s1_translator_avalon_anti_slave_0_clken;                                                  // onchip_memory_0_s1_translator:av_clken -> onchip_memory_0:clken
	wire         onchip_memory_0_s1_translator_avalon_anti_slave_0_write;                                                  // onchip_memory_0_s1_translator:av_write -> onchip_memory_0:write
	wire  [31:0] onchip_memory_0_s1_translator_avalon_anti_slave_0_readdata;                                               // onchip_memory_0:readdata -> onchip_memory_0_s1_translator:av_readdata
	wire   [3:0] onchip_memory_0_s1_translator_avalon_anti_slave_0_byteenable;                                             // onchip_memory_0_s1_translator:av_byteenable -> onchip_memory_0:byteenable
	wire  [31:0] onchip_shared_s1_translator_avalon_anti_slave_0_writedata;                                                // onchip_shared_s1_translator:av_writedata -> onchip_shared:writedata
	wire  [13:0] onchip_shared_s1_translator_avalon_anti_slave_0_address;                                                  // onchip_shared_s1_translator:av_address -> onchip_shared:address
	wire         onchip_shared_s1_translator_avalon_anti_slave_0_chipselect;                                               // onchip_shared_s1_translator:av_chipselect -> onchip_shared:chipselect
	wire         onchip_shared_s1_translator_avalon_anti_slave_0_clken;                                                    // onchip_shared_s1_translator:av_clken -> onchip_shared:clken
	wire         onchip_shared_s1_translator_avalon_anti_slave_0_write;                                                    // onchip_shared_s1_translator:av_write -> onchip_shared:write
	wire  [31:0] onchip_shared_s1_translator_avalon_anti_slave_0_readdata;                                                 // onchip_shared:readdata -> onchip_shared_s1_translator:av_readdata
	wire   [3:0] onchip_shared_s1_translator_avalon_anti_slave_0_byteenable;                                               // onchip_shared_s1_translator:av_byteenable -> onchip_shared:byteenable
	wire  [15:0] timer_0_0_s1_translator_avalon_anti_slave_0_writedata;                                                    // timer_0_0_s1_translator:av_writedata -> timer_0_0:writedata
	wire   [2:0] timer_0_0_s1_translator_avalon_anti_slave_0_address;                                                      // timer_0_0_s1_translator:av_address -> timer_0_0:address
	wire         timer_0_0_s1_translator_avalon_anti_slave_0_chipselect;                                                   // timer_0_0_s1_translator:av_chipselect -> timer_0_0:chipselect
	wire         timer_0_0_s1_translator_avalon_anti_slave_0_write;                                                        // timer_0_0_s1_translator:av_write -> timer_0_0:write_n
	wire  [15:0] timer_0_0_s1_translator_avalon_anti_slave_0_readdata;                                                     // timer_0_0:readdata -> timer_0_0_s1_translator:av_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                 // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                   // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                     // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                  // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                       // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                        // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                    // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire  [31:0] mutex_0_s1_translator_avalon_anti_slave_0_writedata;                                                      // mutex_0_s1_translator:av_writedata -> mutex_0:data_from_cpu
	wire   [0:0] mutex_0_s1_translator_avalon_anti_slave_0_address;                                                        // mutex_0_s1_translator:av_address -> mutex_0:address
	wire         mutex_0_s1_translator_avalon_anti_slave_0_chipselect;                                                     // mutex_0_s1_translator:av_chipselect -> mutex_0:chipselect
	wire         mutex_0_s1_translator_avalon_anti_slave_0_write;                                                          // mutex_0_s1_translator:av_write -> mutex_0:write
	wire         mutex_0_s1_translator_avalon_anti_slave_0_read;                                                           // mutex_0_s1_translator:av_read -> mutex_0:read
	wire  [31:0] mutex_0_s1_translator_avalon_anti_slave_0_readdata;                                                       // mutex_0:data_to_cpu -> mutex_0_s1_translator:av_readdata
	wire  [31:0] mutex_1_s1_translator_avalon_anti_slave_0_writedata;                                                      // mutex_1_s1_translator:av_writedata -> mutex_1:data_from_cpu
	wire   [0:0] mutex_1_s1_translator_avalon_anti_slave_0_address;                                                        // mutex_1_s1_translator:av_address -> mutex_1:address
	wire         mutex_1_s1_translator_avalon_anti_slave_0_chipselect;                                                     // mutex_1_s1_translator:av_chipselect -> mutex_1:chipselect
	wire         mutex_1_s1_translator_avalon_anti_slave_0_write;                                                          // mutex_1_s1_translator:av_write -> mutex_1:write
	wire         mutex_1_s1_translator_avalon_anti_slave_0_read;                                                           // mutex_1_s1_translator:av_read -> mutex_1:read
	wire  [31:0] mutex_1_s1_translator_avalon_anti_slave_0_readdata;                                                       // mutex_1:data_to_cpu -> mutex_1_s1_translator:av_readdata
	wire  [31:0] mutex_2_s1_translator_avalon_anti_slave_0_writedata;                                                      // mutex_2_s1_translator:av_writedata -> mutex_2:data_from_cpu
	wire   [0:0] mutex_2_s1_translator_avalon_anti_slave_0_address;                                                        // mutex_2_s1_translator:av_address -> mutex_2:address
	wire         mutex_2_s1_translator_avalon_anti_slave_0_chipselect;                                                     // mutex_2_s1_translator:av_chipselect -> mutex_2:chipselect
	wire         mutex_2_s1_translator_avalon_anti_slave_0_write;                                                          // mutex_2_s1_translator:av_write -> mutex_2:write
	wire         mutex_2_s1_translator_avalon_anti_slave_0_read;                                                           // mutex_2_s1_translator:av_read -> mutex_2:read
	wire  [31:0] mutex_2_s1_translator_avalon_anti_slave_0_readdata;                                                       // mutex_2:data_to_cpu -> mutex_2_s1_translator:av_readdata
	wire  [31:0] mutex_3_s1_translator_avalon_anti_slave_0_writedata;                                                      // mutex_3_s1_translator:av_writedata -> mutex_3:data_from_cpu
	wire   [0:0] mutex_3_s1_translator_avalon_anti_slave_0_address;                                                        // mutex_3_s1_translator:av_address -> mutex_3:address
	wire         mutex_3_s1_translator_avalon_anti_slave_0_chipselect;                                                     // mutex_3_s1_translator:av_chipselect -> mutex_3:chipselect
	wire         mutex_3_s1_translator_avalon_anti_slave_0_write;                                                          // mutex_3_s1_translator:av_write -> mutex_3:write
	wire         mutex_3_s1_translator_avalon_anti_slave_0_read;                                                           // mutex_3_s1_translator:av_read -> mutex_3:read
	wire  [31:0] mutex_3_s1_translator_avalon_anti_slave_0_readdata;                                                       // mutex_3:data_to_cpu -> mutex_3_s1_translator:av_readdata
	wire  [31:0] mutex_4_s1_translator_avalon_anti_slave_0_writedata;                                                      // mutex_4_s1_translator:av_writedata -> mutex_4:data_from_cpu
	wire   [0:0] mutex_4_s1_translator_avalon_anti_slave_0_address;                                                        // mutex_4_s1_translator:av_address -> mutex_4:address
	wire         mutex_4_s1_translator_avalon_anti_slave_0_chipselect;                                                     // mutex_4_s1_translator:av_chipselect -> mutex_4:chipselect
	wire         mutex_4_s1_translator_avalon_anti_slave_0_write;                                                          // mutex_4_s1_translator:av_write -> mutex_4:write
	wire         mutex_4_s1_translator_avalon_anti_slave_0_read;                                                           // mutex_4_s1_translator:av_read -> mutex_4:read
	wire  [31:0] mutex_4_s1_translator_avalon_anti_slave_0_readdata;                                                       // mutex_4:data_to_cpu -> mutex_4_s1_translator:av_readdata
	wire  [31:0] mutex_5_s1_translator_avalon_anti_slave_0_writedata;                                                      // mutex_5_s1_translator:av_writedata -> mutex_5:data_from_cpu
	wire   [0:0] mutex_5_s1_translator_avalon_anti_slave_0_address;                                                        // mutex_5_s1_translator:av_address -> mutex_5:address
	wire         mutex_5_s1_translator_avalon_anti_slave_0_chipselect;                                                     // mutex_5_s1_translator:av_chipselect -> mutex_5:chipselect
	wire         mutex_5_s1_translator_avalon_anti_slave_0_write;                                                          // mutex_5_s1_translator:av_write -> mutex_5:write
	wire         mutex_5_s1_translator_avalon_anti_slave_0_read;                                                           // mutex_5_s1_translator:av_read -> mutex_5:read
	wire  [31:0] mutex_5_s1_translator_avalon_anti_slave_0_readdata;                                                       // mutex_5:data_to_cpu -> mutex_5_s1_translator:av_readdata
	wire         fifo_0_to_1_in_translator_avalon_anti_slave_0_waitrequest;                                                // fifo_0_to_1:avalonmm_write_slave_waitrequest -> fifo_0_to_1_in_translator:av_waitrequest
	wire  [31:0] fifo_0_to_1_in_translator_avalon_anti_slave_0_writedata;                                                  // fifo_0_to_1_in_translator:av_writedata -> fifo_0_to_1:avalonmm_write_slave_writedata
	wire         fifo_0_to_1_in_translator_avalon_anti_slave_0_write;                                                      // fifo_0_to_1_in_translator:av_write -> fifo_0_to_1:avalonmm_write_slave_write
	wire  [31:0] fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_writedata;                                              // fifo_0_to_1_in_csr_translator:av_writedata -> fifo_0_to_1:wrclk_control_slave_writedata
	wire   [2:0] fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_address;                                                // fifo_0_to_1_in_csr_translator:av_address -> fifo_0_to_1:wrclk_control_slave_address
	wire         fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_write;                                                  // fifo_0_to_1_in_csr_translator:av_write -> fifo_0_to_1:wrclk_control_slave_write
	wire         fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_read;                                                   // fifo_0_to_1_in_csr_translator:av_read -> fifo_0_to_1:wrclk_control_slave_read
	wire  [31:0] fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_readdata;                                               // fifo_0_to_1:wrclk_control_slave_readdata -> fifo_0_to_1_in_csr_translator:av_readdata
	wire         fifo_0_to_2_in_translator_avalon_anti_slave_0_waitrequest;                                                // fifo_0_to_2:avalonmm_write_slave_waitrequest -> fifo_0_to_2_in_translator:av_waitrequest
	wire  [31:0] fifo_0_to_2_in_translator_avalon_anti_slave_0_writedata;                                                  // fifo_0_to_2_in_translator:av_writedata -> fifo_0_to_2:avalonmm_write_slave_writedata
	wire         fifo_0_to_2_in_translator_avalon_anti_slave_0_write;                                                      // fifo_0_to_2_in_translator:av_write -> fifo_0_to_2:avalonmm_write_slave_write
	wire  [31:0] fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_writedata;                                              // fifo_0_to_2_in_csr_translator:av_writedata -> fifo_0_to_2:wrclk_control_slave_writedata
	wire   [2:0] fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_address;                                                // fifo_0_to_2_in_csr_translator:av_address -> fifo_0_to_2:wrclk_control_slave_address
	wire         fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_write;                                                  // fifo_0_to_2_in_csr_translator:av_write -> fifo_0_to_2:wrclk_control_slave_write
	wire         fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_read;                                                   // fifo_0_to_2_in_csr_translator:av_read -> fifo_0_to_2:wrclk_control_slave_read
	wire  [31:0] fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_readdata;                                               // fifo_0_to_2:wrclk_control_slave_readdata -> fifo_0_to_2_in_csr_translator:av_readdata
	wire  [31:0] fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_writedata;                                             // fifo_1_to_0_out_csr_translator:av_writedata -> fifo_1_to_0:rdclk_control_slave_writedata
	wire   [2:0] fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_address;                                               // fifo_1_to_0_out_csr_translator:av_address -> fifo_1_to_0:rdclk_control_slave_address
	wire         fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_write;                                                 // fifo_1_to_0_out_csr_translator:av_write -> fifo_1_to_0:rdclk_control_slave_write
	wire         fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_read;                                                  // fifo_1_to_0_out_csr_translator:av_read -> fifo_1_to_0:rdclk_control_slave_read
	wire  [31:0] fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_readdata;                                              // fifo_1_to_0:rdclk_control_slave_readdata -> fifo_1_to_0_out_csr_translator:av_readdata
	wire         fifo_1_to_0_out_translator_avalon_anti_slave_0_waitrequest;                                               // fifo_1_to_0:avalonmm_read_slave_waitrequest -> fifo_1_to_0_out_translator:av_waitrequest
	wire         fifo_1_to_0_out_translator_avalon_anti_slave_0_read;                                                      // fifo_1_to_0_out_translator:av_read -> fifo_1_to_0:avalonmm_read_slave_read
	wire  [31:0] fifo_1_to_0_out_translator_avalon_anti_slave_0_readdata;                                                  // fifo_1_to_0:avalonmm_read_slave_readdata -> fifo_1_to_0_out_translator:av_readdata
	wire         fifo_2_to_0_out_translator_avalon_anti_slave_0_waitrequest;                                               // fifo_2_to_0:avalonmm_read_slave_waitrequest -> fifo_2_to_0_out_translator:av_waitrequest
	wire         fifo_2_to_0_out_translator_avalon_anti_slave_0_read;                                                      // fifo_2_to_0_out_translator:av_read -> fifo_2_to_0:avalonmm_read_slave_read
	wire  [31:0] fifo_2_to_0_out_translator_avalon_anti_slave_0_readdata;                                                  // fifo_2_to_0:avalonmm_read_slave_readdata -> fifo_2_to_0_out_translator:av_readdata
	wire  [31:0] fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_writedata;                                             // fifo_2_to_0_out_csr_translator:av_writedata -> fifo_2_to_0:rdclk_control_slave_writedata
	wire   [2:0] fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_address;                                               // fifo_2_to_0_out_csr_translator:av_address -> fifo_2_to_0:rdclk_control_slave_address
	wire         fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_write;                                                 // fifo_2_to_0_out_csr_translator:av_write -> fifo_2_to_0:rdclk_control_slave_write
	wire         fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_read;                                                  // fifo_2_to_0_out_csr_translator:av_read -> fifo_2_to_0:rdclk_control_slave_read
	wire  [31:0] fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_readdata;                                              // fifo_2_to_0:rdclk_control_slave_readdata -> fifo_2_to_0_out_csr_translator:av_readdata
	wire  [31:0] red_leds_s1_translator_avalon_anti_slave_0_writedata;                                                     // red_leds_s1_translator:av_writedata -> red_leds:writedata
	wire   [1:0] red_leds_s1_translator_avalon_anti_slave_0_address;                                                       // red_leds_s1_translator:av_address -> red_leds:address
	wire         red_leds_s1_translator_avalon_anti_slave_0_chipselect;                                                    // red_leds_s1_translator:av_chipselect -> red_leds:chipselect
	wire         red_leds_s1_translator_avalon_anti_slave_0_write;                                                         // red_leds_s1_translator:av_write -> red_leds:write_n
	wire  [31:0] red_leds_s1_translator_avalon_anti_slave_0_readdata;                                                      // red_leds:readdata -> red_leds_s1_translator:av_readdata
	wire  [31:0] green_leds_s1_translator_avalon_anti_slave_0_writedata;                                                   // green_leds_s1_translator:av_writedata -> green_leds:writedata
	wire   [1:0] green_leds_s1_translator_avalon_anti_slave_0_address;                                                     // green_leds_s1_translator:av_address -> green_leds:address
	wire         green_leds_s1_translator_avalon_anti_slave_0_chipselect;                                                  // green_leds_s1_translator:av_chipselect -> green_leds:chipselect
	wire         green_leds_s1_translator_avalon_anti_slave_0_write;                                                       // green_leds_s1_translator:av_write -> green_leds:write_n
	wire  [31:0] green_leds_s1_translator_avalon_anti_slave_0_readdata;                                                    // green_leds:readdata -> green_leds_s1_translator:av_readdata
	wire   [1:0] switches_s1_translator_avalon_anti_slave_0_address;                                                       // switches_s1_translator:av_address -> switches:address
	wire  [31:0] switches_s1_translator_avalon_anti_slave_0_readdata;                                                      // switches:readdata -> switches_s1_translator:av_readdata
	wire  [15:0] timer_shared_0_s1_translator_avalon_anti_slave_0_writedata;                                               // timer_shared_0_s1_translator:av_writedata -> timer_shared_0:writedata
	wire   [2:0] timer_shared_0_s1_translator_avalon_anti_slave_0_address;                                                 // timer_shared_0_s1_translator:av_address -> timer_shared_0:address
	wire         timer_shared_0_s1_translator_avalon_anti_slave_0_chipselect;                                              // timer_shared_0_s1_translator:av_chipselect -> timer_shared_0:chipselect
	wire         timer_shared_0_s1_translator_avalon_anti_slave_0_write;                                                   // timer_shared_0_s1_translator:av_write -> timer_shared_0:write_n
	wire  [15:0] timer_shared_0_s1_translator_avalon_anti_slave_0_readdata;                                                // timer_shared_0:readdata -> timer_shared_0_s1_translator:av_readdata
	wire  [31:0] performance_counter_0_control_slave_translator_avalon_anti_slave_0_writedata;                             // performance_counter_0_control_slave_translator:av_writedata -> performance_counter_0:writedata
	wire   [4:0] performance_counter_0_control_slave_translator_avalon_anti_slave_0_address;                               // performance_counter_0_control_slave_translator:av_address -> performance_counter_0:address
	wire         performance_counter_0_control_slave_translator_avalon_anti_slave_0_write;                                 // performance_counter_0_control_slave_translator:av_write -> performance_counter_0:write
	wire  [31:0] performance_counter_0_control_slave_translator_avalon_anti_slave_0_readdata;                              // performance_counter_0:readdata -> performance_counter_0_control_slave_translator:av_readdata
	wire         performance_counter_0_control_slave_translator_avalon_anti_slave_0_begintransfer;                         // performance_counter_0_control_slave_translator:av_begintransfer -> performance_counter_0:begintransfer
	wire  [15:0] timer_0_1_s1_translator_avalon_anti_slave_0_writedata;                                                    // timer_0_1_s1_translator:av_writedata -> timer_0_1:writedata
	wire   [2:0] timer_0_1_s1_translator_avalon_anti_slave_0_address;                                                      // timer_0_1_s1_translator:av_address -> timer_0_1:address
	wire         timer_0_1_s1_translator_avalon_anti_slave_0_chipselect;                                                   // timer_0_1_s1_translator:av_chipselect -> timer_0_1:chipselect
	wire         timer_0_1_s1_translator_avalon_anti_slave_0_write;                                                        // timer_0_1_s1_translator:av_write -> timer_0_1:write_n
	wire  [15:0] timer_0_1_s1_translator_avalon_anti_slave_0_readdata;                                                     // timer_0_1:readdata -> timer_0_1_s1_translator:av_readdata
	wire  [15:0] timer_shared_1_s1_translator_avalon_anti_slave_0_writedata;                                               // timer_shared_1_s1_translator:av_writedata -> timer_shared_1:writedata
	wire   [2:0] timer_shared_1_s1_translator_avalon_anti_slave_0_address;                                                 // timer_shared_1_s1_translator:av_address -> timer_shared_1:address
	wire         timer_shared_1_s1_translator_avalon_anti_slave_0_chipselect;                                              // timer_shared_1_s1_translator:av_chipselect -> timer_shared_1:chipselect
	wire         timer_shared_1_s1_translator_avalon_anti_slave_0_write;                                                   // timer_shared_1_s1_translator:av_write -> timer_shared_1:write_n
	wire  [15:0] timer_shared_1_s1_translator_avalon_anti_slave_0_readdata;                                                // timer_shared_1:readdata -> timer_shared_1_s1_translator:av_readdata
	wire         cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                       // cpu_1:jtag_debug_module_waitrequest -> cpu_1_jtag_debug_module_translator:av_waitrequest
	wire  [31:0] cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                         // cpu_1_jtag_debug_module_translator:av_writedata -> cpu_1:jtag_debug_module_writedata
	wire   [8:0] cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_address;                                           // cpu_1_jtag_debug_module_translator:av_address -> cpu_1:jtag_debug_module_address
	wire         cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_write;                                             // cpu_1_jtag_debug_module_translator:av_write -> cpu_1:jtag_debug_module_write
	wire         cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_read;                                              // cpu_1_jtag_debug_module_translator:av_read -> cpu_1:jtag_debug_module_read
	wire  [31:0] cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                          // cpu_1:jtag_debug_module_readdata -> cpu_1_jtag_debug_module_translator:av_readdata
	wire         cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                       // cpu_1_jtag_debug_module_translator:av_debugaccess -> cpu_1:jtag_debug_module_debugaccess
	wire   [3:0] cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                        // cpu_1_jtag_debug_module_translator:av_byteenable -> cpu_1:jtag_debug_module_byteenable
	wire  [31:0] onchip_memory_1_s1_translator_avalon_anti_slave_0_writedata;                                              // onchip_memory_1_s1_translator:av_writedata -> onchip_memory_1:writedata
	wire  [12:0] onchip_memory_1_s1_translator_avalon_anti_slave_0_address;                                                // onchip_memory_1_s1_translator:av_address -> onchip_memory_1:address
	wire         onchip_memory_1_s1_translator_avalon_anti_slave_0_chipselect;                                             // onchip_memory_1_s1_translator:av_chipselect -> onchip_memory_1:chipselect
	wire         onchip_memory_1_s1_translator_avalon_anti_slave_0_clken;                                                  // onchip_memory_1_s1_translator:av_clken -> onchip_memory_1:clken
	wire         onchip_memory_1_s1_translator_avalon_anti_slave_0_write;                                                  // onchip_memory_1_s1_translator:av_write -> onchip_memory_1:write
	wire  [31:0] onchip_memory_1_s1_translator_avalon_anti_slave_0_readdata;                                               // onchip_memory_1:readdata -> onchip_memory_1_s1_translator:av_readdata
	wire   [3:0] onchip_memory_1_s1_translator_avalon_anti_slave_0_byteenable;                                             // onchip_memory_1_s1_translator:av_byteenable -> onchip_memory_1:byteenable
	wire  [15:0] timer_1_0_s1_translator_avalon_anti_slave_0_writedata;                                                    // timer_1_0_s1_translator:av_writedata -> timer_1_0:writedata
	wire   [2:0] timer_1_0_s1_translator_avalon_anti_slave_0_address;                                                      // timer_1_0_s1_translator:av_address -> timer_1_0:address
	wire         timer_1_0_s1_translator_avalon_anti_slave_0_chipselect;                                                   // timer_1_0_s1_translator:av_chipselect -> timer_1_0:chipselect
	wire         timer_1_0_s1_translator_avalon_anti_slave_0_write;                                                        // timer_1_0_s1_translator:av_write -> timer_1_0:write_n
	wire  [15:0] timer_1_0_s1_translator_avalon_anti_slave_0_readdata;                                                     // timer_1_0:readdata -> timer_1_0_s1_translator:av_readdata
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                 // jtag_uart_1:av_waitrequest -> jtag_uart_1_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                   // jtag_uart_1_avalon_jtag_slave_translator:av_writedata -> jtag_uart_1:av_writedata
	wire   [0:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                     // jtag_uart_1_avalon_jtag_slave_translator:av_address -> jtag_uart_1:av_address
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                  // jtag_uart_1_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_1:av_chipselect
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                       // jtag_uart_1_avalon_jtag_slave_translator:av_write -> jtag_uart_1:av_write_n
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                        // jtag_uart_1_avalon_jtag_slave_translator:av_read -> jtag_uart_1:av_read_n
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                    // jtag_uart_1:av_readdata -> jtag_uart_1_avalon_jtag_slave_translator:av_readdata
	wire         fifo_0_to_1_out_translator_avalon_anti_slave_0_waitrequest;                                               // fifo_0_to_1:avalonmm_read_slave_waitrequest -> fifo_0_to_1_out_translator:av_waitrequest
	wire         fifo_0_to_1_out_translator_avalon_anti_slave_0_read;                                                      // fifo_0_to_1_out_translator:av_read -> fifo_0_to_1:avalonmm_read_slave_read
	wire  [31:0] fifo_0_to_1_out_translator_avalon_anti_slave_0_readdata;                                                  // fifo_0_to_1:avalonmm_read_slave_readdata -> fifo_0_to_1_out_translator:av_readdata
	wire  [31:0] fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_writedata;                                             // fifo_0_to_1_out_csr_translator:av_writedata -> fifo_0_to_1:rdclk_control_slave_writedata
	wire   [2:0] fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_address;                                               // fifo_0_to_1_out_csr_translator:av_address -> fifo_0_to_1:rdclk_control_slave_address
	wire         fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_write;                                                 // fifo_0_to_1_out_csr_translator:av_write -> fifo_0_to_1:rdclk_control_slave_write
	wire         fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_read;                                                  // fifo_0_to_1_out_csr_translator:av_read -> fifo_0_to_1:rdclk_control_slave_read
	wire  [31:0] fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_readdata;                                              // fifo_0_to_1:rdclk_control_slave_readdata -> fifo_0_to_1_out_csr_translator:av_readdata
	wire         fifo_1_to_0_in_translator_avalon_anti_slave_0_waitrequest;                                                // fifo_1_to_0:avalonmm_write_slave_waitrequest -> fifo_1_to_0_in_translator:av_waitrequest
	wire  [31:0] fifo_1_to_0_in_translator_avalon_anti_slave_0_writedata;                                                  // fifo_1_to_0_in_translator:av_writedata -> fifo_1_to_0:avalonmm_write_slave_writedata
	wire         fifo_1_to_0_in_translator_avalon_anti_slave_0_write;                                                      // fifo_1_to_0_in_translator:av_write -> fifo_1_to_0:avalonmm_write_slave_write
	wire  [31:0] fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_writedata;                                              // fifo_1_to_0_in_csr_translator:av_writedata -> fifo_1_to_0:wrclk_control_slave_writedata
	wire   [2:0] fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_address;                                                // fifo_1_to_0_in_csr_translator:av_address -> fifo_1_to_0:wrclk_control_slave_address
	wire         fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_write;                                                  // fifo_1_to_0_in_csr_translator:av_write -> fifo_1_to_0:wrclk_control_slave_write
	wire         fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_read;                                                   // fifo_1_to_0_in_csr_translator:av_read -> fifo_1_to_0:wrclk_control_slave_read
	wire  [31:0] fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_readdata;                                               // fifo_1_to_0:wrclk_control_slave_readdata -> fifo_1_to_0_in_csr_translator:av_readdata
	wire         fifo_1_to_2_in_translator_avalon_anti_slave_0_waitrequest;                                                // fifo_1_to_2:avalonmm_write_slave_waitrequest -> fifo_1_to_2_in_translator:av_waitrequest
	wire  [31:0] fifo_1_to_2_in_translator_avalon_anti_slave_0_writedata;                                                  // fifo_1_to_2_in_translator:av_writedata -> fifo_1_to_2:avalonmm_write_slave_writedata
	wire         fifo_1_to_2_in_translator_avalon_anti_slave_0_write;                                                      // fifo_1_to_2_in_translator:av_write -> fifo_1_to_2:avalonmm_write_slave_write
	wire  [31:0] fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_writedata;                                              // fifo_1_to_2_in_csr_translator:av_writedata -> fifo_1_to_2:wrclk_control_slave_writedata
	wire   [2:0] fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_address;                                                // fifo_1_to_2_in_csr_translator:av_address -> fifo_1_to_2:wrclk_control_slave_address
	wire         fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_write;                                                  // fifo_1_to_2_in_csr_translator:av_write -> fifo_1_to_2:wrclk_control_slave_write
	wire         fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_read;                                                   // fifo_1_to_2_in_csr_translator:av_read -> fifo_1_to_2:wrclk_control_slave_read
	wire  [31:0] fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_readdata;                                               // fifo_1_to_2:wrclk_control_slave_readdata -> fifo_1_to_2_in_csr_translator:av_readdata
	wire         fifo_2_to_1_out_translator_avalon_anti_slave_0_waitrequest;                                               // fifo_2_to_1:avalonmm_read_slave_waitrequest -> fifo_2_to_1_out_translator:av_waitrequest
	wire         fifo_2_to_1_out_translator_avalon_anti_slave_0_read;                                                      // fifo_2_to_1_out_translator:av_read -> fifo_2_to_1:avalonmm_read_slave_read
	wire  [31:0] fifo_2_to_1_out_translator_avalon_anti_slave_0_readdata;                                                  // fifo_2_to_1:avalonmm_read_slave_readdata -> fifo_2_to_1_out_translator:av_readdata
	wire  [31:0] fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_writedata;                                             // fifo_2_to_1_out_csr_translator:av_writedata -> fifo_2_to_1:rdclk_control_slave_writedata
	wire   [2:0] fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_address;                                               // fifo_2_to_1_out_csr_translator:av_address -> fifo_2_to_1:rdclk_control_slave_address
	wire         fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_write;                                                 // fifo_2_to_1_out_csr_translator:av_write -> fifo_2_to_1:rdclk_control_slave_write
	wire         fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_read;                                                  // fifo_2_to_1_out_csr_translator:av_read -> fifo_2_to_1:rdclk_control_slave_read
	wire  [31:0] fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_readdata;                                              // fifo_2_to_1:rdclk_control_slave_readdata -> fifo_2_to_1_out_csr_translator:av_readdata
	wire  [31:0] performance_counter_1_control_slave_translator_avalon_anti_slave_0_writedata;                             // performance_counter_1_control_slave_translator:av_writedata -> performance_counter_1:writedata
	wire   [4:0] performance_counter_1_control_slave_translator_avalon_anti_slave_0_address;                               // performance_counter_1_control_slave_translator:av_address -> performance_counter_1:address
	wire         performance_counter_1_control_slave_translator_avalon_anti_slave_0_write;                                 // performance_counter_1_control_slave_translator:av_write -> performance_counter_1:write
	wire  [31:0] performance_counter_1_control_slave_translator_avalon_anti_slave_0_readdata;                              // performance_counter_1:readdata -> performance_counter_1_control_slave_translator:av_readdata
	wire         performance_counter_1_control_slave_translator_avalon_anti_slave_0_begintransfer;                         // performance_counter_1_control_slave_translator:av_begintransfer -> performance_counter_1:begintransfer
	wire  [15:0] timer_1_1_s1_translator_avalon_anti_slave_0_writedata;                                                    // timer_1_1_s1_translator:av_writedata -> timer_1_1:writedata
	wire   [2:0] timer_1_1_s1_translator_avalon_anti_slave_0_address;                                                      // timer_1_1_s1_translator:av_address -> timer_1_1:address
	wire         timer_1_1_s1_translator_avalon_anti_slave_0_chipselect;                                                   // timer_1_1_s1_translator:av_chipselect -> timer_1_1:chipselect
	wire         timer_1_1_s1_translator_avalon_anti_slave_0_write;                                                        // timer_1_1_s1_translator:av_write -> timer_1_1:write_n
	wire  [15:0] timer_1_1_s1_translator_avalon_anti_slave_0_readdata;                                                     // timer_1_1:readdata -> timer_1_1_s1_translator:av_readdata
	wire         cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                       // cpu_2:jtag_debug_module_waitrequest -> cpu_2_jtag_debug_module_translator:av_waitrequest
	wire  [31:0] cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                         // cpu_2_jtag_debug_module_translator:av_writedata -> cpu_2:jtag_debug_module_writedata
	wire   [8:0] cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_address;                                           // cpu_2_jtag_debug_module_translator:av_address -> cpu_2:jtag_debug_module_address
	wire         cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_write;                                             // cpu_2_jtag_debug_module_translator:av_write -> cpu_2:jtag_debug_module_write
	wire         cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_read;                                              // cpu_2_jtag_debug_module_translator:av_read -> cpu_2:jtag_debug_module_read
	wire  [31:0] cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                          // cpu_2:jtag_debug_module_readdata -> cpu_2_jtag_debug_module_translator:av_readdata
	wire         cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                       // cpu_2_jtag_debug_module_translator:av_debugaccess -> cpu_2:jtag_debug_module_debugaccess
	wire   [3:0] cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                        // cpu_2_jtag_debug_module_translator:av_byteenable -> cpu_2:jtag_debug_module_byteenable
	wire  [31:0] onchip_memory_2_s1_translator_avalon_anti_slave_0_writedata;                                              // onchip_memory_2_s1_translator:av_writedata -> onchip_memory_2:writedata
	wire  [12:0] onchip_memory_2_s1_translator_avalon_anti_slave_0_address;                                                // onchip_memory_2_s1_translator:av_address -> onchip_memory_2:address
	wire         onchip_memory_2_s1_translator_avalon_anti_slave_0_chipselect;                                             // onchip_memory_2_s1_translator:av_chipselect -> onchip_memory_2:chipselect
	wire         onchip_memory_2_s1_translator_avalon_anti_slave_0_clken;                                                  // onchip_memory_2_s1_translator:av_clken -> onchip_memory_2:clken
	wire         onchip_memory_2_s1_translator_avalon_anti_slave_0_write;                                                  // onchip_memory_2_s1_translator:av_write -> onchip_memory_2:write
	wire  [31:0] onchip_memory_2_s1_translator_avalon_anti_slave_0_readdata;                                               // onchip_memory_2:readdata -> onchip_memory_2_s1_translator:av_readdata
	wire   [3:0] onchip_memory_2_s1_translator_avalon_anti_slave_0_byteenable;                                             // onchip_memory_2_s1_translator:av_byteenable -> onchip_memory_2:byteenable
	wire  [15:0] timer_2_0_s1_translator_avalon_anti_slave_0_writedata;                                                    // timer_2_0_s1_translator:av_writedata -> timer_2_0:writedata
	wire   [2:0] timer_2_0_s1_translator_avalon_anti_slave_0_address;                                                      // timer_2_0_s1_translator:av_address -> timer_2_0:address
	wire         timer_2_0_s1_translator_avalon_anti_slave_0_chipselect;                                                   // timer_2_0_s1_translator:av_chipselect -> timer_2_0:chipselect
	wire         timer_2_0_s1_translator_avalon_anti_slave_0_write;                                                        // timer_2_0_s1_translator:av_write -> timer_2_0:write_n
	wire  [15:0] timer_2_0_s1_translator_avalon_anti_slave_0_readdata;                                                     // timer_2_0:readdata -> timer_2_0_s1_translator:av_readdata
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                 // jtag_uart_2:av_waitrequest -> jtag_uart_2_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                   // jtag_uart_2_avalon_jtag_slave_translator:av_writedata -> jtag_uart_2:av_writedata
	wire   [0:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                     // jtag_uart_2_avalon_jtag_slave_translator:av_address -> jtag_uart_2:av_address
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                  // jtag_uart_2_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_2:av_chipselect
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                       // jtag_uart_2_avalon_jtag_slave_translator:av_write -> jtag_uart_2:av_write_n
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                        // jtag_uart_2_avalon_jtag_slave_translator:av_read -> jtag_uart_2:av_read_n
	wire  [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                    // jtag_uart_2:av_readdata -> jtag_uart_2_avalon_jtag_slave_translator:av_readdata
	wire         fifo_0_to_2_out_translator_avalon_anti_slave_0_waitrequest;                                               // fifo_0_to_2:avalonmm_read_slave_waitrequest -> fifo_0_to_2_out_translator:av_waitrequest
	wire         fifo_0_to_2_out_translator_avalon_anti_slave_0_read;                                                      // fifo_0_to_2_out_translator:av_read -> fifo_0_to_2:avalonmm_read_slave_read
	wire  [31:0] fifo_0_to_2_out_translator_avalon_anti_slave_0_readdata;                                                  // fifo_0_to_2:avalonmm_read_slave_readdata -> fifo_0_to_2_out_translator:av_readdata
	wire  [31:0] fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_writedata;                                             // fifo_0_to_2_out_csr_translator:av_writedata -> fifo_0_to_2:rdclk_control_slave_writedata
	wire   [2:0] fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_address;                                               // fifo_0_to_2_out_csr_translator:av_address -> fifo_0_to_2:rdclk_control_slave_address
	wire         fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_write;                                                 // fifo_0_to_2_out_csr_translator:av_write -> fifo_0_to_2:rdclk_control_slave_write
	wire         fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_read;                                                  // fifo_0_to_2_out_csr_translator:av_read -> fifo_0_to_2:rdclk_control_slave_read
	wire  [31:0] fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_readdata;                                              // fifo_0_to_2:rdclk_control_slave_readdata -> fifo_0_to_2_out_csr_translator:av_readdata
	wire         fifo_1_to_2_out_translator_avalon_anti_slave_0_waitrequest;                                               // fifo_1_to_2:avalonmm_read_slave_waitrequest -> fifo_1_to_2_out_translator:av_waitrequest
	wire         fifo_1_to_2_out_translator_avalon_anti_slave_0_read;                                                      // fifo_1_to_2_out_translator:av_read -> fifo_1_to_2:avalonmm_read_slave_read
	wire  [31:0] fifo_1_to_2_out_translator_avalon_anti_slave_0_readdata;                                                  // fifo_1_to_2:avalonmm_read_slave_readdata -> fifo_1_to_2_out_translator:av_readdata
	wire  [31:0] fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_writedata;                                             // fifo_1_to_2_out_csr_translator:av_writedata -> fifo_1_to_2:rdclk_control_slave_writedata
	wire   [2:0] fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_address;                                               // fifo_1_to_2_out_csr_translator:av_address -> fifo_1_to_2:rdclk_control_slave_address
	wire         fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_write;                                                 // fifo_1_to_2_out_csr_translator:av_write -> fifo_1_to_2:rdclk_control_slave_write
	wire         fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_read;                                                  // fifo_1_to_2_out_csr_translator:av_read -> fifo_1_to_2:rdclk_control_slave_read
	wire  [31:0] fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_readdata;                                              // fifo_1_to_2:rdclk_control_slave_readdata -> fifo_1_to_2_out_csr_translator:av_readdata
	wire         fifo_2_to_0_in_translator_avalon_anti_slave_0_waitrequest;                                                // fifo_2_to_0:avalonmm_write_slave_waitrequest -> fifo_2_to_0_in_translator:av_waitrequest
	wire  [31:0] fifo_2_to_0_in_translator_avalon_anti_slave_0_writedata;                                                  // fifo_2_to_0_in_translator:av_writedata -> fifo_2_to_0:avalonmm_write_slave_writedata
	wire         fifo_2_to_0_in_translator_avalon_anti_slave_0_write;                                                      // fifo_2_to_0_in_translator:av_write -> fifo_2_to_0:avalonmm_write_slave_write
	wire  [31:0] fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_writedata;                                              // fifo_2_to_0_in_csr_translator:av_writedata -> fifo_2_to_0:wrclk_control_slave_writedata
	wire   [2:0] fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_address;                                                // fifo_2_to_0_in_csr_translator:av_address -> fifo_2_to_0:wrclk_control_slave_address
	wire         fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_write;                                                  // fifo_2_to_0_in_csr_translator:av_write -> fifo_2_to_0:wrclk_control_slave_write
	wire         fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_read;                                                   // fifo_2_to_0_in_csr_translator:av_read -> fifo_2_to_0:wrclk_control_slave_read
	wire  [31:0] fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_readdata;                                               // fifo_2_to_0:wrclk_control_slave_readdata -> fifo_2_to_0_in_csr_translator:av_readdata
	wire         fifo_2_to_1_in_translator_avalon_anti_slave_0_waitrequest;                                                // fifo_2_to_1:avalonmm_write_slave_waitrequest -> fifo_2_to_1_in_translator:av_waitrequest
	wire  [31:0] fifo_2_to_1_in_translator_avalon_anti_slave_0_writedata;                                                  // fifo_2_to_1_in_translator:av_writedata -> fifo_2_to_1:avalonmm_write_slave_writedata
	wire         fifo_2_to_1_in_translator_avalon_anti_slave_0_write;                                                      // fifo_2_to_1_in_translator:av_write -> fifo_2_to_1:avalonmm_write_slave_write
	wire  [31:0] fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_writedata;                                              // fifo_2_to_1_in_csr_translator:av_writedata -> fifo_2_to_1:wrclk_control_slave_writedata
	wire   [2:0] fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_address;                                                // fifo_2_to_1_in_csr_translator:av_address -> fifo_2_to_1:wrclk_control_slave_address
	wire         fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_write;                                                  // fifo_2_to_1_in_csr_translator:av_write -> fifo_2_to_1:wrclk_control_slave_write
	wire         fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_read;                                                   // fifo_2_to_1_in_csr_translator:av_read -> fifo_2_to_1:wrclk_control_slave_read
	wire  [31:0] fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_readdata;                                               // fifo_2_to_1:wrclk_control_slave_readdata -> fifo_2_to_1_in_csr_translator:av_readdata
	wire  [31:0] performance_counter_2_control_slave_translator_avalon_anti_slave_0_writedata;                             // performance_counter_2_control_slave_translator:av_writedata -> performance_counter_2:writedata
	wire   [4:0] performance_counter_2_control_slave_translator_avalon_anti_slave_0_address;                               // performance_counter_2_control_slave_translator:av_address -> performance_counter_2:address
	wire         performance_counter_2_control_slave_translator_avalon_anti_slave_0_write;                                 // performance_counter_2_control_slave_translator:av_write -> performance_counter_2:write
	wire  [31:0] performance_counter_2_control_slave_translator_avalon_anti_slave_0_readdata;                              // performance_counter_2:readdata -> performance_counter_2_control_slave_translator:av_readdata
	wire         performance_counter_2_control_slave_translator_avalon_anti_slave_0_begintransfer;                         // performance_counter_2_control_slave_translator:av_begintransfer -> performance_counter_2:begintransfer
	wire  [15:0] timer_2_1_s1_translator_avalon_anti_slave_0_writedata;                                                    // timer_2_1_s1_translator:av_writedata -> timer_2_1:writedata
	wire   [2:0] timer_2_1_s1_translator_avalon_anti_slave_0_address;                                                      // timer_2_1_s1_translator:av_address -> timer_2_1:address
	wire         timer_2_1_s1_translator_avalon_anti_slave_0_chipselect;                                                   // timer_2_1_s1_translator:av_chipselect -> timer_2_1:chipselect
	wire         timer_2_1_s1_translator_avalon_anti_slave_0_write;                                                        // timer_2_1_s1_translator:av_write -> timer_2_1:write_n
	wire  [15:0] timer_2_1_s1_translator_avalon_anti_slave_0_readdata;                                                     // timer_2_1:readdata -> timer_2_1_s1_translator:av_readdata
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                                // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount;                                 // cpu_0_instruction_master_translator:uav_burstcount -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_writedata;                                  // cpu_0_instruction_master_translator:uav_writedata -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [17:0] cpu_0_instruction_master_translator_avalon_universal_master_0_address;                                    // cpu_0_instruction_master_translator:uav_address -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_lock;                                       // cpu_0_instruction_master_translator:uav_lock -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_write;                                      // cpu_0_instruction_master_translator:uav_write -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_read;                                       // cpu_0_instruction_master_translator:uav_read -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_readdata;                                   // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_instruction_master_translator:uav_readdata
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                                // cpu_0_instruction_master_translator:uav_debugaccess -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable;                                 // cpu_0_instruction_master_translator:uav_byteenable -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                              // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_instruction_master_translator:uav_readdatavalid
	wire         cpu_0_data_master_translator_avalon_universal_master_0_waitrequest;                                       // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_0_data_master_translator_avalon_universal_master_0_burstcount;                                        // cpu_0_data_master_translator:uav_burstcount -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_0_data_master_translator_avalon_universal_master_0_writedata;                                         // cpu_0_data_master_translator:uav_writedata -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [17:0] cpu_0_data_master_translator_avalon_universal_master_0_address;                                           // cpu_0_data_master_translator:uav_address -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_0_data_master_translator_avalon_universal_master_0_lock;                                              // cpu_0_data_master_translator:uav_lock -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_0_data_master_translator_avalon_universal_master_0_write;                                             // cpu_0_data_master_translator:uav_write -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_0_data_master_translator_avalon_universal_master_0_read;                                              // cpu_0_data_master_translator:uav_read -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_0_data_master_translator_avalon_universal_master_0_readdata;                                          // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_data_master_translator:uav_readdata
	wire         cpu_0_data_master_translator_avalon_universal_master_0_debugaccess;                                       // cpu_0_data_master_translator:uav_debugaccess -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_0_data_master_translator_avalon_universal_master_0_byteenable;                                        // cpu_0_data_master_translator:uav_byteenable -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid;                                     // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_data_master_translator:uav_readdatavalid
	wire         cpu_1_data_master_translator_avalon_universal_master_0_waitrequest;                                       // cpu_1_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_1_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_1_data_master_translator_avalon_universal_master_0_burstcount;                                        // cpu_1_data_master_translator:uav_burstcount -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_1_data_master_translator_avalon_universal_master_0_writedata;                                         // cpu_1_data_master_translator:uav_writedata -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [17:0] cpu_1_data_master_translator_avalon_universal_master_0_address;                                           // cpu_1_data_master_translator:uav_address -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_1_data_master_translator_avalon_universal_master_0_lock;                                              // cpu_1_data_master_translator:uav_lock -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_1_data_master_translator_avalon_universal_master_0_write;                                             // cpu_1_data_master_translator:uav_write -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_1_data_master_translator_avalon_universal_master_0_read;                                              // cpu_1_data_master_translator:uav_read -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_1_data_master_translator_avalon_universal_master_0_readdata;                                          // cpu_1_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_1_data_master_translator:uav_readdata
	wire         cpu_1_data_master_translator_avalon_universal_master_0_debugaccess;                                       // cpu_1_data_master_translator:uav_debugaccess -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_1_data_master_translator_avalon_universal_master_0_byteenable;                                        // cpu_1_data_master_translator:uav_byteenable -> cpu_1_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_1_data_master_translator_avalon_universal_master_0_readdatavalid;                                     // cpu_1_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_1_data_master_translator:uav_readdatavalid
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_waitrequest;                                // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_1_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_1_instruction_master_translator_avalon_universal_master_0_burstcount;                                 // cpu_1_instruction_master_translator:uav_burstcount -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_1_instruction_master_translator_avalon_universal_master_0_writedata;                                  // cpu_1_instruction_master_translator:uav_writedata -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [17:0] cpu_1_instruction_master_translator_avalon_universal_master_0_address;                                    // cpu_1_instruction_master_translator:uav_address -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_lock;                                       // cpu_1_instruction_master_translator:uav_lock -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_write;                                      // cpu_1_instruction_master_translator:uav_write -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_read;                                       // cpu_1_instruction_master_translator:uav_read -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_1_instruction_master_translator_avalon_universal_master_0_readdata;                                   // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_1_instruction_master_translator:uav_readdata
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_debugaccess;                                // cpu_1_instruction_master_translator:uav_debugaccess -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_1_instruction_master_translator_avalon_universal_master_0_byteenable;                                 // cpu_1_instruction_master_translator:uav_byteenable -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_readdatavalid;                              // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_1_instruction_master_translator:uav_readdatavalid
	wire         cpu_2_data_master_translator_avalon_universal_master_0_waitrequest;                                       // cpu_2_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_2_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_2_data_master_translator_avalon_universal_master_0_burstcount;                                        // cpu_2_data_master_translator:uav_burstcount -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_2_data_master_translator_avalon_universal_master_0_writedata;                                         // cpu_2_data_master_translator:uav_writedata -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [17:0] cpu_2_data_master_translator_avalon_universal_master_0_address;                                           // cpu_2_data_master_translator:uav_address -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_2_data_master_translator_avalon_universal_master_0_lock;                                              // cpu_2_data_master_translator:uav_lock -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_2_data_master_translator_avalon_universal_master_0_write;                                             // cpu_2_data_master_translator:uav_write -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_2_data_master_translator_avalon_universal_master_0_read;                                              // cpu_2_data_master_translator:uav_read -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_2_data_master_translator_avalon_universal_master_0_readdata;                                          // cpu_2_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_2_data_master_translator:uav_readdata
	wire         cpu_2_data_master_translator_avalon_universal_master_0_debugaccess;                                       // cpu_2_data_master_translator:uav_debugaccess -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_2_data_master_translator_avalon_universal_master_0_byteenable;                                        // cpu_2_data_master_translator:uav_byteenable -> cpu_2_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_2_data_master_translator_avalon_universal_master_0_readdatavalid;                                     // cpu_2_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_2_data_master_translator:uav_readdatavalid
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_waitrequest;                                // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_2_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_2_instruction_master_translator_avalon_universal_master_0_burstcount;                                 // cpu_2_instruction_master_translator:uav_burstcount -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_2_instruction_master_translator_avalon_universal_master_0_writedata;                                  // cpu_2_instruction_master_translator:uav_writedata -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [17:0] cpu_2_instruction_master_translator_avalon_universal_master_0_address;                                    // cpu_2_instruction_master_translator:uav_address -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_lock;                                       // cpu_2_instruction_master_translator:uav_lock -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_write;                                      // cpu_2_instruction_master_translator:uav_write -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_read;                                       // cpu_2_instruction_master_translator:uav_read -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_2_instruction_master_translator_avalon_universal_master_0_readdata;                                   // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_2_instruction_master_translator:uav_readdata
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_debugaccess;                                // cpu_2_instruction_master_translator:uav_debugaccess -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_2_instruction_master_translator_avalon_universal_master_0_byteenable;                                 // cpu_2_instruction_master_translator:uav_byteenable -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_readdatavalid;                              // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_2_instruction_master_translator:uav_readdatavalid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // cpu_0_jtag_debug_module_translator:uav_waitrequest -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_0_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                           // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_0_jtag_debug_module_translator:uav_writedata
	wire  [17:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                             // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_0_jtag_debug_module_translator:uav_address
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                               // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_0_jtag_debug_module_translator:uav_write
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_0_jtag_debug_module_translator:uav_lock
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_0_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                            // cpu_0_jtag_debug_module_translator:uav_readdata -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // cpu_0_jtag_debug_module_translator:uav_readdatavalid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_0_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_0_jtag_debug_module_translator:uav_byteenable
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                         // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // onchip_memory_0_s1_translator:uav_waitrequest -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory_0_s1_translator:uav_burstcount
	wire  [31:0] onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory_0_s1_translator:uav_writedata
	wire  [17:0] onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory_0_s1_translator:uav_address
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory_0_s1_translator:uav_write
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory_0_s1_translator:uav_lock
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory_0_s1_translator:uav_read
	wire  [31:0] onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // onchip_memory_0_s1_translator:uav_readdata -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // onchip_memory_0_s1_translator:uav_readdatavalid -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory_0_s1_translator:uav_debugaccess
	wire   [3:0] onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory_0_s1_translator:uav_byteenable
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // onchip_shared_s1_translator:uav_waitrequest -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // onchip_shared_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_shared_s1_translator:uav_burstcount
	wire  [31:0] onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // onchip_shared_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_shared_s1_translator:uav_writedata
	wire  [17:0] onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // onchip_shared_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_shared_s1_translator:uav_address
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // onchip_shared_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_shared_s1_translator:uav_write
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // onchip_shared_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_shared_s1_translator:uav_lock
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // onchip_shared_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_shared_s1_translator:uav_read
	wire  [31:0] onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // onchip_shared_s1_translator:uav_readdata -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // onchip_shared_s1_translator:uav_readdatavalid -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // onchip_shared_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_shared_s1_translator:uav_debugaccess
	wire   [3:0] onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // onchip_shared_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_shared_s1_translator:uav_byteenable
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // onchip_shared_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // onchip_shared_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // onchip_shared_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // onchip_shared_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // onchip_shared_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // onchip_shared_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] onchip_shared_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // onchip_shared_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // onchip_shared_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // timer_0_0_s1_translator:uav_waitrequest -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // timer_0_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_0_s1_translator:uav_burstcount
	wire  [31:0] timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // timer_0_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_0_s1_translator:uav_writedata
	wire  [17:0] timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // timer_0_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_0_s1_translator:uav_address
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // timer_0_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_0_s1_translator:uav_write
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // timer_0_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_0_s1_translator:uav_lock
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // timer_0_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_0_s1_translator:uav_read
	wire  [31:0] timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // timer_0_0_s1_translator:uav_readdata -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // timer_0_0_s1_translator:uav_readdatavalid -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // timer_0_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // timer_0_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_0_s1_translator:uav_byteenable
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // timer_0_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // timer_0_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // timer_0_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // timer_0_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // timer_0_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // timer_0_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_0_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // timer_0_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // timer_0_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire  [17:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                      // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // mutex_0_s1_translator:uav_waitrequest -> mutex_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // mutex_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> mutex_0_s1_translator:uav_burstcount
	wire  [31:0] mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // mutex_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> mutex_0_s1_translator:uav_writedata
	wire  [17:0] mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // mutex_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> mutex_0_s1_translator:uav_address
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // mutex_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> mutex_0_s1_translator:uav_write
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // mutex_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> mutex_0_s1_translator:uav_lock
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // mutex_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> mutex_0_s1_translator:uav_read
	wire  [31:0] mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // mutex_0_s1_translator:uav_readdata -> mutex_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // mutex_0_s1_translator:uav_readdatavalid -> mutex_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // mutex_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mutex_0_s1_translator:uav_debugaccess
	wire   [3:0] mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // mutex_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> mutex_0_s1_translator:uav_byteenable
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // mutex_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // mutex_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // mutex_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // mutex_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mutex_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mutex_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mutex_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mutex_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mutex_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // mutex_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // mutex_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mutex_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] mutex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // mutex_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mutex_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // mutex_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mutex_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // mutex_1_s1_translator:uav_waitrequest -> mutex_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // mutex_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> mutex_1_s1_translator:uav_burstcount
	wire  [31:0] mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // mutex_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> mutex_1_s1_translator:uav_writedata
	wire  [17:0] mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // mutex_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> mutex_1_s1_translator:uav_address
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // mutex_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> mutex_1_s1_translator:uav_write
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // mutex_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> mutex_1_s1_translator:uav_lock
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // mutex_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> mutex_1_s1_translator:uav_read
	wire  [31:0] mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // mutex_1_s1_translator:uav_readdata -> mutex_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // mutex_1_s1_translator:uav_readdatavalid -> mutex_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // mutex_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mutex_1_s1_translator:uav_debugaccess
	wire   [3:0] mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // mutex_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> mutex_1_s1_translator:uav_byteenable
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // mutex_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // mutex_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // mutex_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // mutex_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mutex_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mutex_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mutex_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mutex_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mutex_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // mutex_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // mutex_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mutex_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] mutex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // mutex_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mutex_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // mutex_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mutex_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // mutex_2_s1_translator:uav_waitrequest -> mutex_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // mutex_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> mutex_2_s1_translator:uav_burstcount
	wire  [31:0] mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // mutex_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> mutex_2_s1_translator:uav_writedata
	wire  [17:0] mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // mutex_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> mutex_2_s1_translator:uav_address
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // mutex_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> mutex_2_s1_translator:uav_write
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // mutex_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> mutex_2_s1_translator:uav_lock
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // mutex_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> mutex_2_s1_translator:uav_read
	wire  [31:0] mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // mutex_2_s1_translator:uav_readdata -> mutex_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // mutex_2_s1_translator:uav_readdatavalid -> mutex_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // mutex_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mutex_2_s1_translator:uav_debugaccess
	wire   [3:0] mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // mutex_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> mutex_2_s1_translator:uav_byteenable
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // mutex_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // mutex_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // mutex_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // mutex_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mutex_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mutex_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mutex_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mutex_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mutex_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // mutex_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // mutex_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mutex_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] mutex_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // mutex_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mutex_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // mutex_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mutex_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // mutex_3_s1_translator:uav_waitrequest -> mutex_3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // mutex_3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> mutex_3_s1_translator:uav_burstcount
	wire  [31:0] mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // mutex_3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> mutex_3_s1_translator:uav_writedata
	wire  [17:0] mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // mutex_3_s1_translator_avalon_universal_slave_0_agent:m0_address -> mutex_3_s1_translator:uav_address
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // mutex_3_s1_translator_avalon_universal_slave_0_agent:m0_write -> mutex_3_s1_translator:uav_write
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // mutex_3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> mutex_3_s1_translator:uav_lock
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // mutex_3_s1_translator_avalon_universal_slave_0_agent:m0_read -> mutex_3_s1_translator:uav_read
	wire  [31:0] mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // mutex_3_s1_translator:uav_readdata -> mutex_3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // mutex_3_s1_translator:uav_readdatavalid -> mutex_3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // mutex_3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mutex_3_s1_translator:uav_debugaccess
	wire   [3:0] mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // mutex_3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> mutex_3_s1_translator:uav_byteenable
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // mutex_3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // mutex_3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // mutex_3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // mutex_3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mutex_3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mutex_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mutex_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mutex_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mutex_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // mutex_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // mutex_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mutex_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] mutex_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // mutex_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mutex_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // mutex_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mutex_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // mutex_4_s1_translator:uav_waitrequest -> mutex_4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // mutex_4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> mutex_4_s1_translator:uav_burstcount
	wire  [31:0] mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // mutex_4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> mutex_4_s1_translator:uav_writedata
	wire  [17:0] mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // mutex_4_s1_translator_avalon_universal_slave_0_agent:m0_address -> mutex_4_s1_translator:uav_address
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // mutex_4_s1_translator_avalon_universal_slave_0_agent:m0_write -> mutex_4_s1_translator:uav_write
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // mutex_4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> mutex_4_s1_translator:uav_lock
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // mutex_4_s1_translator_avalon_universal_slave_0_agent:m0_read -> mutex_4_s1_translator:uav_read
	wire  [31:0] mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // mutex_4_s1_translator:uav_readdata -> mutex_4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // mutex_4_s1_translator:uav_readdatavalid -> mutex_4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // mutex_4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mutex_4_s1_translator:uav_debugaccess
	wire   [3:0] mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // mutex_4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> mutex_4_s1_translator:uav_byteenable
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // mutex_4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // mutex_4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // mutex_4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // mutex_4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mutex_4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mutex_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mutex_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mutex_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mutex_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // mutex_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // mutex_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mutex_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] mutex_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // mutex_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mutex_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // mutex_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mutex_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // mutex_5_s1_translator:uav_waitrequest -> mutex_5_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // mutex_5_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> mutex_5_s1_translator:uav_burstcount
	wire  [31:0] mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // mutex_5_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> mutex_5_s1_translator:uav_writedata
	wire  [17:0] mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // mutex_5_s1_translator_avalon_universal_slave_0_agent:m0_address -> mutex_5_s1_translator:uav_address
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // mutex_5_s1_translator_avalon_universal_slave_0_agent:m0_write -> mutex_5_s1_translator:uav_write
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // mutex_5_s1_translator_avalon_universal_slave_0_agent:m0_lock -> mutex_5_s1_translator:uav_lock
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // mutex_5_s1_translator_avalon_universal_slave_0_agent:m0_read -> mutex_5_s1_translator:uav_read
	wire  [31:0] mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // mutex_5_s1_translator:uav_readdata -> mutex_5_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // mutex_5_s1_translator:uav_readdatavalid -> mutex_5_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // mutex_5_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mutex_5_s1_translator:uav_debugaccess
	wire   [3:0] mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // mutex_5_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> mutex_5_s1_translator:uav_byteenable
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // mutex_5_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // mutex_5_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // mutex_5_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // mutex_5_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mutex_5_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mutex_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mutex_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mutex_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mutex_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // mutex_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // mutex_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mutex_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] mutex_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // mutex_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mutex_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // mutex_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mutex_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // fifo_0_to_1_in_translator:uav_waitrequest -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_to_1_in_translator:uav_burstcount
	wire  [31:0] fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_to_1_in_translator:uav_writedata
	wire  [17:0] fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_address;                                      // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_to_1_in_translator:uav_address
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_write;                                        // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_to_1_in_translator:uav_write
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_lock;                                         // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_to_1_in_translator:uav_lock
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_read;                                         // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_to_1_in_translator:uav_read
	wire  [31:0] fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // fifo_0_to_1_in_translator:uav_readdata -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // fifo_0_to_1_in_translator:uav_readdatavalid -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_to_1_in_translator:uav_debugaccess
	wire   [3:0] fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_to_1_in_translator:uav_byteenable
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // fifo_0_to_1_in_csr_translator:uav_waitrequest -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_to_1_in_csr_translator:uav_burstcount
	wire  [31:0] fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_to_1_in_csr_translator:uav_writedata
	wire  [17:0] fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                  // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_to_1_in_csr_translator:uav_address
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                    // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_to_1_in_csr_translator:uav_write
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                     // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_to_1_in_csr_translator:uav_lock
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                     // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_to_1_in_csr_translator:uav_read
	wire  [31:0] fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // fifo_0_to_1_in_csr_translator:uav_readdata -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // fifo_0_to_1_in_csr_translator:uav_readdatavalid -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_to_1_in_csr_translator:uav_debugaccess
	wire   [3:0] fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_to_1_in_csr_translator:uav_byteenable
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                              // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // fifo_0_to_2_in_translator:uav_waitrequest -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_to_2_in_translator:uav_burstcount
	wire  [31:0] fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_to_2_in_translator:uav_writedata
	wire  [17:0] fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_address;                                      // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_to_2_in_translator:uav_address
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_write;                                        // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_to_2_in_translator:uav_write
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock;                                         // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_to_2_in_translator:uav_lock
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_read;                                         // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_to_2_in_translator:uav_read
	wire  [31:0] fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // fifo_0_to_2_in_translator:uav_readdata -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // fifo_0_to_2_in_translator:uav_readdatavalid -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_to_2_in_translator:uav_debugaccess
	wire   [3:0] fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_to_2_in_translator:uav_byteenable
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // fifo_0_to_2_in_csr_translator:uav_waitrequest -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_to_2_in_csr_translator:uav_burstcount
	wire  [31:0] fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_to_2_in_csr_translator:uav_writedata
	wire  [17:0] fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                  // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_to_2_in_csr_translator:uav_address
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                    // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_to_2_in_csr_translator:uav_write
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                     // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_to_2_in_csr_translator:uav_lock
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                     // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_to_2_in_csr_translator:uav_read
	wire  [31:0] fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // fifo_0_to_2_in_csr_translator:uav_readdata -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // fifo_0_to_2_in_csr_translator:uav_readdatavalid -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_to_2_in_csr_translator:uav_debugaccess
	wire   [3:0] fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_to_2_in_csr_translator:uav_byteenable
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                              // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // fifo_1_to_0_out_csr_translator:uav_waitrequest -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_1_to_0_out_csr_translator:uav_burstcount
	wire  [31:0] fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_1_to_0_out_csr_translator:uav_writedata
	wire  [17:0] fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_1_to_0_out_csr_translator:uav_address
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_1_to_0_out_csr_translator:uav_write
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_1_to_0_out_csr_translator:uav_lock
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_1_to_0_out_csr_translator:uav_read
	wire  [31:0] fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // fifo_1_to_0_out_csr_translator:uav_readdata -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // fifo_1_to_0_out_csr_translator:uav_readdatavalid -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_1_to_0_out_csr_translator:uav_debugaccess
	wire   [3:0] fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_1_to_0_out_csr_translator:uav_byteenable
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // fifo_1_to_0_out_translator:uav_waitrequest -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_1_to_0_out_translator:uav_burstcount
	wire  [31:0] fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_1_to_0_out_translator:uav_writedata
	wire  [17:0] fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_address;                                     // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_1_to_0_out_translator:uav_address
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_write;                                       // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_1_to_0_out_translator:uav_write
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_lock;                                        // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_1_to_0_out_translator:uav_lock
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_read;                                        // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_1_to_0_out_translator:uav_read
	wire  [31:0] fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // fifo_1_to_0_out_translator:uav_readdata -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // fifo_1_to_0_out_translator:uav_readdatavalid -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_1_to_0_out_translator:uav_debugaccess
	wire   [3:0] fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_1_to_0_out_translator:uav_byteenable
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // fifo_2_to_0_out_translator:uav_waitrequest -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_2_to_0_out_translator:uav_burstcount
	wire  [31:0] fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_2_to_0_out_translator:uav_writedata
	wire  [17:0] fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_address;                                     // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_2_to_0_out_translator:uav_address
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_write;                                       // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_2_to_0_out_translator:uav_write
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_lock;                                        // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_2_to_0_out_translator:uav_lock
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_read;                                        // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_2_to_0_out_translator:uav_read
	wire  [31:0] fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // fifo_2_to_0_out_translator:uav_readdata -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // fifo_2_to_0_out_translator:uav_readdatavalid -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_2_to_0_out_translator:uav_debugaccess
	wire   [3:0] fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_2_to_0_out_translator:uav_byteenable
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // fifo_2_to_0_out_csr_translator:uav_waitrequest -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_2_to_0_out_csr_translator:uav_burstcount
	wire  [31:0] fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_2_to_0_out_csr_translator:uav_writedata
	wire  [17:0] fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_2_to_0_out_csr_translator:uav_address
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_2_to_0_out_csr_translator:uav_write
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_2_to_0_out_csr_translator:uav_lock
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_2_to_0_out_csr_translator:uav_read
	wire  [31:0] fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // fifo_2_to_0_out_csr_translator:uav_readdata -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // fifo_2_to_0_out_csr_translator:uav_readdatavalid -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_2_to_0_out_csr_translator:uav_debugaccess
	wire   [3:0] fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_2_to_0_out_csr_translator:uav_byteenable
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // red_leds_s1_translator:uav_waitrequest -> red_leds_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] red_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> red_leds_s1_translator:uav_burstcount
	wire  [31:0] red_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> red_leds_s1_translator:uav_writedata
	wire  [17:0] red_leds_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_address -> red_leds_s1_translator:uav_address
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_write -> red_leds_s1_translator:uav_write
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_lock -> red_leds_s1_translator:uav_lock
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_read -> red_leds_s1_translator:uav_read
	wire  [31:0] red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // red_leds_s1_translator:uav_readdata -> red_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // red_leds_s1_translator:uav_readdatavalid -> red_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> red_leds_s1_translator:uav_debugaccess
	wire   [3:0] red_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // red_leds_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> red_leds_s1_translator:uav_byteenable
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // green_leds_s1_translator:uav_waitrequest -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> green_leds_s1_translator:uav_burstcount
	wire  [31:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> green_leds_s1_translator:uav_writedata
	wire  [17:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_address -> green_leds_s1_translator:uav_address
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_write -> green_leds_s1_translator:uav_write
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_lock -> green_leds_s1_translator:uav_lock
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_read -> green_leds_s1_translator:uav_read
	wire  [31:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // green_leds_s1_translator:uav_readdata -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // green_leds_s1_translator:uav_readdatavalid -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> green_leds_s1_translator:uav_debugaccess
	wire   [3:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> green_leds_s1_translator:uav_byteenable
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // switches_s1_translator:uav_waitrequest -> switches_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // switches_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switches_s1_translator:uav_burstcount
	wire  [31:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // switches_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switches_s1_translator:uav_writedata
	wire  [17:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // switches_s1_translator_avalon_universal_slave_0_agent:m0_address -> switches_s1_translator:uav_address
	wire         switches_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // switches_s1_translator_avalon_universal_slave_0_agent:m0_write -> switches_s1_translator:uav_write
	wire         switches_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // switches_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switches_s1_translator:uav_lock
	wire         switches_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // switches_s1_translator_avalon_universal_slave_0_agent:m0_read -> switches_s1_translator:uav_read
	wire  [31:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // switches_s1_translator:uav_readdata -> switches_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // switches_s1_translator:uav_readdatavalid -> switches_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // switches_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switches_s1_translator:uav_debugaccess
	wire   [3:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // switches_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switches_s1_translator:uav_byteenable
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // switches_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // switches_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // switches_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // switches_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switches_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // timer_shared_0_s1_translator:uav_waitrequest -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_shared_0_s1_translator:uav_burstcount
	wire  [31:0] timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_shared_0_s1_translator:uav_writedata
	wire  [17:0] timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_shared_0_s1_translator:uav_address
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_shared_0_s1_translator:uav_write
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_shared_0_s1_translator:uav_lock
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_shared_0_s1_translator:uav_read
	wire  [31:0] timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // timer_shared_0_s1_translator:uav_readdata -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // timer_shared_0_s1_translator:uav_readdatavalid -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_shared_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_shared_0_s1_translator:uav_byteenable
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // performance_counter_0_control_slave_translator:uav_waitrequest -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> performance_counter_0_control_slave_translator:uav_burstcount
	wire  [31:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> performance_counter_0_control_slave_translator:uav_writedata
	wire  [17:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> performance_counter_0_control_slave_translator:uav_address
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> performance_counter_0_control_slave_translator:uav_write
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> performance_counter_0_control_slave_translator:uav_lock
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> performance_counter_0_control_slave_translator:uav_read
	wire  [31:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // performance_counter_0_control_slave_translator:uav_readdata -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // performance_counter_0_control_slave_translator:uav_readdatavalid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> performance_counter_0_control_slave_translator:uav_debugaccess
	wire   [3:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> performance_counter_0_control_slave_translator:uav_byteenable
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // timer_0_1_s1_translator:uav_waitrequest -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // timer_0_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_1_s1_translator:uav_burstcount
	wire  [31:0] timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // timer_0_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_1_s1_translator:uav_writedata
	wire  [17:0] timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // timer_0_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_1_s1_translator:uav_address
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // timer_0_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_1_s1_translator:uav_write
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // timer_0_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_1_s1_translator:uav_lock
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // timer_0_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_1_s1_translator:uav_read
	wire  [31:0] timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // timer_0_1_s1_translator:uav_readdata -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // timer_0_1_s1_translator:uav_readdatavalid -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // timer_0_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_1_s1_translator:uav_debugaccess
	wire   [3:0] timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // timer_0_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_1_s1_translator:uav_byteenable
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // timer_0_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // timer_0_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // timer_0_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // timer_0_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // timer_0_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // timer_0_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_0_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // timer_0_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // timer_0_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // timer_shared_1_s1_translator:uav_waitrequest -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_shared_1_s1_translator:uav_burstcount
	wire  [31:0] timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_shared_1_s1_translator:uav_writedata
	wire  [17:0] timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_shared_1_s1_translator:uav_address
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_shared_1_s1_translator:uav_write
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_shared_1_s1_translator:uav_lock
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_shared_1_s1_translator:uav_read
	wire  [31:0] timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // timer_shared_1_s1_translator:uav_readdata -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // timer_shared_1_s1_translator:uav_readdatavalid -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_shared_1_s1_translator:uav_debugaccess
	wire   [3:0] timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_shared_1_s1_translator:uav_byteenable
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // cpu_1_jtag_debug_module_translator:uav_waitrequest -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_1_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                           // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_1_jtag_debug_module_translator:uav_writedata
	wire  [17:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                             // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_1_jtag_debug_module_translator:uav_address
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                               // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_1_jtag_debug_module_translator:uav_write
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_1_jtag_debug_module_translator:uav_lock
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_1_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                            // cpu_1_jtag_debug_module_translator:uav_readdata -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // cpu_1_jtag_debug_module_translator:uav_readdatavalid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_1_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_1_jtag_debug_module_translator:uav_byteenable
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                         // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // onchip_memory_1_s1_translator:uav_waitrequest -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory_1_s1_translator:uav_burstcount
	wire  [31:0] onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory_1_s1_translator:uav_writedata
	wire  [17:0] onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory_1_s1_translator:uav_address
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory_1_s1_translator:uav_write
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory_1_s1_translator:uav_lock
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory_1_s1_translator:uav_read
	wire  [31:0] onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // onchip_memory_1_s1_translator:uav_readdata -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // onchip_memory_1_s1_translator:uav_readdatavalid -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory_1_s1_translator:uav_debugaccess
	wire   [3:0] onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory_1_s1_translator:uav_byteenable
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // timer_1_0_s1_translator:uav_waitrequest -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // timer_1_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_1_0_s1_translator:uav_burstcount
	wire  [31:0] timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // timer_1_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_1_0_s1_translator:uav_writedata
	wire  [17:0] timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // timer_1_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_1_0_s1_translator:uav_address
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // timer_1_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_1_0_s1_translator:uav_write
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // timer_1_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_1_0_s1_translator:uav_lock
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // timer_1_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_1_0_s1_translator:uav_read
	wire  [31:0] timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // timer_1_0_s1_translator:uav_readdata -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // timer_1_0_s1_translator:uav_readdatavalid -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // timer_1_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_1_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // timer_1_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_1_0_s1_translator:uav_byteenable
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // timer_1_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // timer_1_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // timer_1_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // timer_1_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // timer_1_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // timer_1_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_1_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // timer_1_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // timer_1_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // jtag_uart_1_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_1_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                     // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_1_avalon_jtag_slave_translator:uav_writedata
	wire  [17:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                       // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_1_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                         // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_1_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                          // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_1_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                          // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_1_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                      // jtag_uart_1_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // jtag_uart_1_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_1_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_1_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                   // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // fifo_0_to_1_out_translator:uav_waitrequest -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_to_1_out_translator:uav_burstcount
	wire  [31:0] fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_to_1_out_translator:uav_writedata
	wire  [17:0] fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_address;                                     // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_to_1_out_translator:uav_address
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_write;                                       // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_to_1_out_translator:uav_write
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_lock;                                        // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_to_1_out_translator:uav_lock
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_read;                                        // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_to_1_out_translator:uav_read
	wire  [31:0] fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // fifo_0_to_1_out_translator:uav_readdata -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // fifo_0_to_1_out_translator:uav_readdatavalid -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_to_1_out_translator:uav_debugaccess
	wire   [3:0] fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_to_1_out_translator:uav_byteenable
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // fifo_0_to_1_out_csr_translator:uav_waitrequest -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_to_1_out_csr_translator:uav_burstcount
	wire  [31:0] fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_to_1_out_csr_translator:uav_writedata
	wire  [17:0] fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_to_1_out_csr_translator:uav_address
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_to_1_out_csr_translator:uav_write
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_to_1_out_csr_translator:uav_lock
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_to_1_out_csr_translator:uav_read
	wire  [31:0] fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // fifo_0_to_1_out_csr_translator:uav_readdata -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // fifo_0_to_1_out_csr_translator:uav_readdatavalid -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_to_1_out_csr_translator:uav_debugaccess
	wire   [3:0] fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_to_1_out_csr_translator:uav_byteenable
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // fifo_1_to_0_in_translator:uav_waitrequest -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_1_to_0_in_translator:uav_burstcount
	wire  [31:0] fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_1_to_0_in_translator:uav_writedata
	wire  [17:0] fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_address;                                      // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_1_to_0_in_translator:uav_address
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_write;                                        // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_1_to_0_in_translator:uav_write
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_lock;                                         // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_1_to_0_in_translator:uav_lock
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_read;                                         // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_1_to_0_in_translator:uav_read
	wire  [31:0] fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // fifo_1_to_0_in_translator:uav_readdata -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // fifo_1_to_0_in_translator:uav_readdatavalid -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_1_to_0_in_translator:uav_debugaccess
	wire   [3:0] fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_1_to_0_in_translator:uav_byteenable
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // fifo_1_to_0_in_csr_translator:uav_waitrequest -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_1_to_0_in_csr_translator:uav_burstcount
	wire  [31:0] fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_1_to_0_in_csr_translator:uav_writedata
	wire  [17:0] fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                  // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_1_to_0_in_csr_translator:uav_address
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                    // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_1_to_0_in_csr_translator:uav_write
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                     // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_1_to_0_in_csr_translator:uav_lock
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                     // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_1_to_0_in_csr_translator:uav_read
	wire  [31:0] fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // fifo_1_to_0_in_csr_translator:uav_readdata -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // fifo_1_to_0_in_csr_translator:uav_readdatavalid -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_1_to_0_in_csr_translator:uav_debugaccess
	wire   [3:0] fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_1_to_0_in_csr_translator:uav_byteenable
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                              // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // fifo_1_to_2_in_translator:uav_waitrequest -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_1_to_2_in_translator:uav_burstcount
	wire  [31:0] fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_1_to_2_in_translator:uav_writedata
	wire  [17:0] fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_address;                                      // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_1_to_2_in_translator:uav_address
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_write;                                        // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_1_to_2_in_translator:uav_write
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock;                                         // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_1_to_2_in_translator:uav_lock
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_read;                                         // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_1_to_2_in_translator:uav_read
	wire  [31:0] fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // fifo_1_to_2_in_translator:uav_readdata -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // fifo_1_to_2_in_translator:uav_readdatavalid -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_1_to_2_in_translator:uav_debugaccess
	wire   [3:0] fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_1_to_2_in_translator:uav_byteenable
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // fifo_1_to_2_in_csr_translator:uav_waitrequest -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_1_to_2_in_csr_translator:uav_burstcount
	wire  [31:0] fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_1_to_2_in_csr_translator:uav_writedata
	wire  [17:0] fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                  // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_1_to_2_in_csr_translator:uav_address
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                    // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_1_to_2_in_csr_translator:uav_write
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                     // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_1_to_2_in_csr_translator:uav_lock
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                     // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_1_to_2_in_csr_translator:uav_read
	wire  [31:0] fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // fifo_1_to_2_in_csr_translator:uav_readdata -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // fifo_1_to_2_in_csr_translator:uav_readdatavalid -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_1_to_2_in_csr_translator:uav_debugaccess
	wire   [3:0] fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_1_to_2_in_csr_translator:uav_byteenable
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                              // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // fifo_2_to_1_out_translator:uav_waitrequest -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_2_to_1_out_translator:uav_burstcount
	wire  [31:0] fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_2_to_1_out_translator:uav_writedata
	wire  [17:0] fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_address;                                     // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_2_to_1_out_translator:uav_address
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_write;                                       // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_2_to_1_out_translator:uav_write
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_lock;                                        // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_2_to_1_out_translator:uav_lock
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_read;                                        // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_2_to_1_out_translator:uav_read
	wire  [31:0] fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // fifo_2_to_1_out_translator:uav_readdata -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // fifo_2_to_1_out_translator:uav_readdatavalid -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_2_to_1_out_translator:uav_debugaccess
	wire   [3:0] fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_2_to_1_out_translator:uav_byteenable
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // fifo_2_to_1_out_csr_translator:uav_waitrequest -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_2_to_1_out_csr_translator:uav_burstcount
	wire  [31:0] fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_2_to_1_out_csr_translator:uav_writedata
	wire  [17:0] fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_2_to_1_out_csr_translator:uav_address
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_2_to_1_out_csr_translator:uav_write
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_2_to_1_out_csr_translator:uav_lock
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_2_to_1_out_csr_translator:uav_read
	wire  [31:0] fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // fifo_2_to_1_out_csr_translator:uav_readdata -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // fifo_2_to_1_out_csr_translator:uav_readdatavalid -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_2_to_1_out_csr_translator:uav_debugaccess
	wire   [3:0] fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_2_to_1_out_csr_translator:uav_byteenable
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // performance_counter_1_control_slave_translator:uav_waitrequest -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> performance_counter_1_control_slave_translator:uav_burstcount
	wire  [31:0] performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> performance_counter_1_control_slave_translator:uav_writedata
	wire  [17:0] performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> performance_counter_1_control_slave_translator:uav_address
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> performance_counter_1_control_slave_translator:uav_write
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> performance_counter_1_control_slave_translator:uav_lock
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> performance_counter_1_control_slave_translator:uav_read
	wire  [31:0] performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // performance_counter_1_control_slave_translator:uav_readdata -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // performance_counter_1_control_slave_translator:uav_readdatavalid -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> performance_counter_1_control_slave_translator:uav_debugaccess
	wire   [3:0] performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> performance_counter_1_control_slave_translator:uav_byteenable
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // timer_1_1_s1_translator:uav_waitrequest -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // timer_1_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_1_1_s1_translator:uav_burstcount
	wire  [31:0] timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // timer_1_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_1_1_s1_translator:uav_writedata
	wire  [17:0] timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // timer_1_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_1_1_s1_translator:uav_address
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // timer_1_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_1_1_s1_translator:uav_write
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // timer_1_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_1_1_s1_translator:uav_lock
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // timer_1_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_1_1_s1_translator:uav_read
	wire  [31:0] timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // timer_1_1_s1_translator:uav_readdata -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // timer_1_1_s1_translator:uav_readdatavalid -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // timer_1_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_1_1_s1_translator:uav_debugaccess
	wire   [3:0] timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // timer_1_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_1_1_s1_translator:uav_byteenable
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // timer_1_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // timer_1_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // timer_1_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // timer_1_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // timer_1_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // timer_1_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_1_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // timer_1_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // timer_1_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // cpu_2_jtag_debug_module_translator:uav_waitrequest -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_2_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                           // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_2_jtag_debug_module_translator:uav_writedata
	wire  [17:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                             // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_2_jtag_debug_module_translator:uav_address
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                               // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_2_jtag_debug_module_translator:uav_write
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_2_jtag_debug_module_translator:uav_lock
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_2_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                            // cpu_2_jtag_debug_module_translator:uav_readdata -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // cpu_2_jtag_debug_module_translator:uav_readdatavalid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_2_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_2_jtag_debug_module_translator:uav_byteenable
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                         // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // onchip_memory_2_s1_translator:uav_waitrequest -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory_2_s1_translator:uav_burstcount
	wire  [31:0] onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory_2_s1_translator:uav_writedata
	wire  [17:0] onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory_2_s1_translator:uav_address
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory_2_s1_translator:uav_write
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory_2_s1_translator:uav_lock
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory_2_s1_translator:uav_read
	wire  [31:0] onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // onchip_memory_2_s1_translator:uav_readdata -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // onchip_memory_2_s1_translator:uav_readdatavalid -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory_2_s1_translator:uav_debugaccess
	wire   [3:0] onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory_2_s1_translator:uav_byteenable
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // timer_2_0_s1_translator:uav_waitrequest -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // timer_2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_2_0_s1_translator:uav_burstcount
	wire  [31:0] timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // timer_2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_2_0_s1_translator:uav_writedata
	wire  [17:0] timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // timer_2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_2_0_s1_translator:uav_address
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // timer_2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_2_0_s1_translator:uav_write
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // timer_2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_2_0_s1_translator:uav_lock
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // timer_2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_2_0_s1_translator:uav_read
	wire  [31:0] timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // timer_2_0_s1_translator:uav_readdata -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // timer_2_0_s1_translator:uav_readdatavalid -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // timer_2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_2_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // timer_2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_2_0_s1_translator:uav_byteenable
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // timer_2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // timer_2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // timer_2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // timer_2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // timer_2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // timer_2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // timer_2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // timer_2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // jtag_uart_2_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_2_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                     // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_2_avalon_jtag_slave_translator:uav_writedata
	wire  [17:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                       // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_2_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                         // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_2_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                          // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_2_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                          // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_2_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                      // jtag_uart_2_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // jtag_uart_2_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_2_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_2_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                   // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // fifo_0_to_2_out_translator:uav_waitrequest -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_to_2_out_translator:uav_burstcount
	wire  [31:0] fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_to_2_out_translator:uav_writedata
	wire  [17:0] fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_address;                                     // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_to_2_out_translator:uav_address
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_write;                                       // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_to_2_out_translator:uav_write
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock;                                        // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_to_2_out_translator:uav_lock
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_read;                                        // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_to_2_out_translator:uav_read
	wire  [31:0] fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // fifo_0_to_2_out_translator:uav_readdata -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // fifo_0_to_2_out_translator:uav_readdatavalid -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_to_2_out_translator:uav_debugaccess
	wire   [3:0] fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_to_2_out_translator:uav_byteenable
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // fifo_0_to_2_out_csr_translator:uav_waitrequest -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_to_2_out_csr_translator:uav_burstcount
	wire  [31:0] fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_to_2_out_csr_translator:uav_writedata
	wire  [17:0] fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_to_2_out_csr_translator:uav_address
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_to_2_out_csr_translator:uav_write
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_to_2_out_csr_translator:uav_lock
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_to_2_out_csr_translator:uav_read
	wire  [31:0] fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // fifo_0_to_2_out_csr_translator:uav_readdata -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // fifo_0_to_2_out_csr_translator:uav_readdatavalid -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_to_2_out_csr_translator:uav_debugaccess
	wire   [3:0] fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_to_2_out_csr_translator:uav_byteenable
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // fifo_1_to_2_out_translator:uav_waitrequest -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_1_to_2_out_translator:uav_burstcount
	wire  [31:0] fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_1_to_2_out_translator:uav_writedata
	wire  [17:0] fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_address;                                     // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:m0_address -> fifo_1_to_2_out_translator:uav_address
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_write;                                       // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:m0_write -> fifo_1_to_2_out_translator:uav_write
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock;                                        // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_1_to_2_out_translator:uav_lock
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_read;                                        // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:m0_read -> fifo_1_to_2_out_translator:uav_read
	wire  [31:0] fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // fifo_1_to_2_out_translator:uav_readdata -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // fifo_1_to_2_out_translator:uav_readdatavalid -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_1_to_2_out_translator:uav_debugaccess
	wire   [3:0] fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_1_to_2_out_translator:uav_byteenable
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // fifo_1_to_2_out_csr_translator:uav_waitrequest -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_1_to_2_out_csr_translator:uav_burstcount
	wire  [31:0] fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_1_to_2_out_csr_translator:uav_writedata
	wire  [17:0] fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_1_to_2_out_csr_translator:uav_address
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_1_to_2_out_csr_translator:uav_write
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_1_to_2_out_csr_translator:uav_lock
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_1_to_2_out_csr_translator:uav_read
	wire  [31:0] fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // fifo_1_to_2_out_csr_translator:uav_readdata -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // fifo_1_to_2_out_csr_translator:uav_readdatavalid -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_1_to_2_out_csr_translator:uav_debugaccess
	wire   [3:0] fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_1_to_2_out_csr_translator:uav_byteenable
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // fifo_2_to_0_in_translator:uav_waitrequest -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_2_to_0_in_translator:uav_burstcount
	wire  [31:0] fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_2_to_0_in_translator:uav_writedata
	wire  [17:0] fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_address;                                      // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_2_to_0_in_translator:uav_address
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_write;                                        // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_2_to_0_in_translator:uav_write
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_lock;                                         // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_2_to_0_in_translator:uav_lock
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_read;                                         // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_2_to_0_in_translator:uav_read
	wire  [31:0] fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // fifo_2_to_0_in_translator:uav_readdata -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // fifo_2_to_0_in_translator:uav_readdatavalid -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_2_to_0_in_translator:uav_debugaccess
	wire   [3:0] fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_2_to_0_in_translator:uav_byteenable
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // fifo_2_to_0_in_csr_translator:uav_waitrequest -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_2_to_0_in_csr_translator:uav_burstcount
	wire  [31:0] fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_2_to_0_in_csr_translator:uav_writedata
	wire  [17:0] fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                  // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_2_to_0_in_csr_translator:uav_address
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                    // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_2_to_0_in_csr_translator:uav_write
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                     // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_2_to_0_in_csr_translator:uav_lock
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                     // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_2_to_0_in_csr_translator:uav_read
	wire  [31:0] fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // fifo_2_to_0_in_csr_translator:uav_readdata -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // fifo_2_to_0_in_csr_translator:uav_readdatavalid -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_2_to_0_in_csr_translator:uav_debugaccess
	wire   [3:0] fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_2_to_0_in_csr_translator:uav_byteenable
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                              // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // fifo_2_to_1_in_translator:uav_waitrequest -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_2_to_1_in_translator:uav_burstcount
	wire  [31:0] fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_2_to_1_in_translator:uav_writedata
	wire  [17:0] fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_address;                                      // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_2_to_1_in_translator:uav_address
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_write;                                        // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_2_to_1_in_translator:uav_write
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_lock;                                         // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_2_to_1_in_translator:uav_lock
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_read;                                         // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_2_to_1_in_translator:uav_read
	wire  [31:0] fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // fifo_2_to_1_in_translator:uav_readdata -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // fifo_2_to_1_in_translator:uav_readdatavalid -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_2_to_1_in_translator:uav_debugaccess
	wire   [3:0] fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_2_to_1_in_translator:uav_byteenable
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // fifo_2_to_1_in_csr_translator:uav_waitrequest -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_2_to_1_in_csr_translator:uav_burstcount
	wire  [31:0] fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_2_to_1_in_csr_translator:uav_writedata
	wire  [17:0] fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                  // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_2_to_1_in_csr_translator:uav_address
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                    // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_2_to_1_in_csr_translator:uav_write
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                     // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_2_to_1_in_csr_translator:uav_lock
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                     // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_2_to_1_in_csr_translator:uav_read
	wire  [31:0] fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // fifo_2_to_1_in_csr_translator:uav_readdata -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // fifo_2_to_1_in_csr_translator:uav_readdatavalid -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_2_to_1_in_csr_translator:uav_debugaccess
	wire   [3:0] fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_2_to_1_in_csr_translator:uav_byteenable
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                              // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // performance_counter_2_control_slave_translator:uav_waitrequest -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> performance_counter_2_control_slave_translator:uav_burstcount
	wire  [31:0] performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> performance_counter_2_control_slave_translator:uav_writedata
	wire  [17:0] performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> performance_counter_2_control_slave_translator:uav_address
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> performance_counter_2_control_slave_translator:uav_write
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> performance_counter_2_control_slave_translator:uav_lock
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> performance_counter_2_control_slave_translator:uav_read
	wire  [31:0] performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // performance_counter_2_control_slave_translator:uav_readdata -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // performance_counter_2_control_slave_translator:uav_readdatavalid -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> performance_counter_2_control_slave_translator:uav_debugaccess
	wire   [3:0] performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> performance_counter_2_control_slave_translator:uav_byteenable
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // timer_2_1_s1_translator:uav_waitrequest -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // timer_2_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_2_1_s1_translator:uav_burstcount
	wire  [31:0] timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // timer_2_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_2_1_s1_translator:uav_writedata
	wire  [17:0] timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // timer_2_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_2_1_s1_translator:uav_address
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // timer_2_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_2_1_s1_translator:uav_write
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // timer_2_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_2_1_s1_translator:uav_lock
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // timer_2_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_2_1_s1_translator:uav_read
	wire  [31:0] timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // timer_2_1_s1_translator:uav_readdata -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // timer_2_1_s1_translator:uav_readdatavalid -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // timer_2_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_2_1_s1_translator:uav_debugaccess
	wire   [3:0] timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // timer_2_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_2_1_s1_translator:uav_byteenable
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // timer_2_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // timer_2_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // timer_2_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [97:0] timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // timer_2_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [97:0] timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // timer_2_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // timer_2_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_2_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // timer_2_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // timer_2_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                             // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [96:0] cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                              // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router:sink_ready -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                              // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                    // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                            // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [96:0] cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                                     // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                    // addr_router_001:sink_ready -> cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                              // cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire         cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                    // cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire         cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                            // cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [96:0] cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_data;                                     // cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire         cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                    // addr_router_002:sink_ready -> cpu_1_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                             // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [96:0] cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                              // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire         cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router_003:sink_ready -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                              // cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire         cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                    // cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire         cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                            // cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [96:0] cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_data;                                     // cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire         cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                    // addr_router_004:sink_ready -> cpu_2_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                             // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire  [96:0] cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                              // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire         cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router_005:sink_ready -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                               // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [96:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router:sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [96:0] onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_001:sink_ready -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // onchip_shared_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // onchip_shared_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // onchip_shared_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [96:0] onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // onchip_shared_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_002:sink_ready -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // timer_0_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // timer_0_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // timer_0_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [96:0] timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // timer_0_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_003:sink_ready -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [96:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_004:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // mutex_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // mutex_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // mutex_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [96:0] mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // mutex_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_005:sink_ready -> mutex_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // mutex_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // mutex_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // mutex_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [96:0] mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // mutex_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_006:sink_ready -> mutex_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // mutex_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // mutex_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // mutex_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [96:0] mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // mutex_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_007:sink_ready -> mutex_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // mutex_3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // mutex_3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // mutex_3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [96:0] mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // mutex_3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_008:sink_ready -> mutex_3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // mutex_4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // mutex_4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // mutex_4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [96:0] mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // mutex_4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_009:sink_ready -> mutex_4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // mutex_5_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // mutex_5_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // mutex_5_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [96:0] mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // mutex_5_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_010:sink_ready -> mutex_5_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_valid;                                        // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [96:0] fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_data;                                         // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire         fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_011:sink_ready -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                    // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [96:0] fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                     // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire         fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_012:sink_ready -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid;                                        // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [96:0] fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_data;                                         // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire         fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_013:sink_ready -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                    // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [96:0] fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                     // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire         fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_014:sink_ready -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [96:0] fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire         fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_015:sink_ready -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_valid;                                       // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [96:0] fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_data;                                        // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire         fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_016:sink_ready -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_valid;                                       // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [96:0] fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_data;                                        // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire         fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_017:sink_ready -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [96:0] fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire         fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_018:sink_ready -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // red_leds_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // red_leds_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // red_leds_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [96:0] red_leds_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // red_leds_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire         red_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_019:sink_ready -> red_leds_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [96:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire         green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_020:sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // switches_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // switches_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // switches_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire  [96:0] switches_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // switches_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire         switches_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_021:sink_ready -> switches_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire  [96:0] timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire         timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_022:sink_ready -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	wire  [96:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	wire         performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_023:sink_ready -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // timer_0_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // timer_0_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // timer_0_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	wire  [96:0] timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // timer_0_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	wire         timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_024:sink_ready -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	wire  [96:0] timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	wire         timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_025:sink_ready -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_026:sink_endofpacket
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                               // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_026:sink_valid
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_026:sink_startofpacket
	wire  [96:0] cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_026:sink_data
	wire         cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_026:sink_ready -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_027:sink_endofpacket
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_027:sink_valid
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_027:sink_startofpacket
	wire  [96:0] onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_027:sink_data
	wire         onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_027:sink_ready -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // timer_1_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_028:sink_endofpacket
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // timer_1_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_028:sink_valid
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // timer_1_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_028:sink_startofpacket
	wire  [96:0] timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // timer_1_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_028:sink_data
	wire         timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_028:sink_ready -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_029:sink_endofpacket
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                         // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_029:sink_valid
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_029:sink_startofpacket
	wire  [96:0] jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                          // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_029:sink_data
	wire         jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_029:sink_ready -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_030:sink_endofpacket
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_valid;                                       // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_030:sink_valid
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_030:sink_startofpacket
	wire  [96:0] fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_data;                                        // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_030:sink_data
	wire         fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_030:sink_ready -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_031:sink_endofpacket
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_031:sink_valid
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_031:sink_startofpacket
	wire  [96:0] fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_031:sink_data
	wire         fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_031:sink_ready -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_032:sink_endofpacket
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_valid;                                        // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_032:sink_valid
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_032:sink_startofpacket
	wire  [96:0] fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_data;                                         // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_032:sink_data
	wire         fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_032:sink_ready -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_033:sink_endofpacket
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                    // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_033:sink_valid
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_033:sink_startofpacket
	wire  [96:0] fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                     // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_033:sink_data
	wire         fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_033:sink_ready -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_034:sink_endofpacket
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid;                                        // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_034:sink_valid
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_034:sink_startofpacket
	wire  [96:0] fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_data;                                         // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_034:sink_data
	wire         fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_034:sink_ready -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_035:sink_endofpacket
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                    // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_035:sink_valid
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_035:sink_startofpacket
	wire  [96:0] fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                     // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_035:sink_data
	wire         fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_035:sink_ready -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_036:sink_endofpacket
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_valid;                                       // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_036:sink_valid
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_036:sink_startofpacket
	wire  [96:0] fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_data;                                        // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_036:sink_data
	wire         fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_036:sink_ready -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_037:sink_endofpacket
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_037:sink_valid
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_037:sink_startofpacket
	wire  [96:0] fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_037:sink_data
	wire         fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_037:sink_ready -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_038:sink_endofpacket
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_038:sink_valid
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_038:sink_startofpacket
	wire  [96:0] performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_038:sink_data
	wire         performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_038:sink_ready -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // timer_1_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_039:sink_endofpacket
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // timer_1_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_039:sink_valid
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // timer_1_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_039:sink_startofpacket
	wire  [96:0] timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // timer_1_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_039:sink_data
	wire         timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_039:sink_ready -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_040:sink_endofpacket
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                               // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_040:sink_valid
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_040:sink_startofpacket
	wire  [96:0] cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_040:sink_data
	wire         cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_040:sink_ready -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_041:sink_endofpacket
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_041:sink_valid
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_041:sink_startofpacket
	wire  [96:0] onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_041:sink_data
	wire         onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_041:sink_ready -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // timer_2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_042:sink_endofpacket
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // timer_2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_042:sink_valid
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // timer_2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_042:sink_startofpacket
	wire  [96:0] timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // timer_2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_042:sink_data
	wire         timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_042:sink_ready -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_043:sink_endofpacket
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                         // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_043:sink_valid
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_043:sink_startofpacket
	wire  [96:0] jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                          // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_043:sink_data
	wire         jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_043:sink_ready -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_044:sink_endofpacket
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid;                                       // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_044:sink_valid
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_044:sink_startofpacket
	wire  [96:0] fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_data;                                        // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_044:sink_data
	wire         fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_044:sink_ready -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_045:sink_endofpacket
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_045:sink_valid
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_045:sink_startofpacket
	wire  [96:0] fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_045:sink_data
	wire         fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_045:sink_ready -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_046:sink_endofpacket
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid;                                       // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_046:sink_valid
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_046:sink_startofpacket
	wire  [96:0] fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_data;                                        // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_046:sink_data
	wire         fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_046:sink_ready -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_047:sink_endofpacket
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_047:sink_valid
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_047:sink_startofpacket
	wire  [96:0] fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_047:sink_data
	wire         fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_047:sink_ready -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_048:sink_endofpacket
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_valid;                                        // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_048:sink_valid
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_048:sink_startofpacket
	wire  [96:0] fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_data;                                         // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_048:sink_data
	wire         fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_048:sink_ready -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_049:sink_endofpacket
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                    // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_049:sink_valid
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_049:sink_startofpacket
	wire  [96:0] fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                     // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_049:sink_data
	wire         fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_049:sink_ready -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_050:sink_endofpacket
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_valid;                                        // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_050:sink_valid
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_050:sink_startofpacket
	wire  [96:0] fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_data;                                         // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_050:sink_data
	wire         fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_050:sink_ready -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_051:sink_endofpacket
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                    // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_051:sink_valid
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_051:sink_startofpacket
	wire  [96:0] fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                     // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_051:sink_data
	wire         fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_051:sink_ready -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_052:sink_endofpacket
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_052:sink_valid
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_052:sink_startofpacket
	wire  [96:0] performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_052:sink_data
	wire         performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_052:sink_ready -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // timer_2_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_053:sink_endofpacket
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // timer_2_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_053:sink_valid
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // timer_2_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_053:sink_startofpacket
	wire  [96:0] timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // timer_2_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_053:sink_data
	wire         timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_053:sink_ready -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rst_controller_reset_out_reset;                                                                           // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cpu_0:reset_n, cpu_0_data_master_translator:reset, cpu_0_data_master_translator_avalon_universal_master_0_agent:reset, cpu_0_instruction_master_translator:reset, cpu_0_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_0_jtag_debug_module_translator:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_0_to_1:wrreset_n, fifo_0_to_1_in_csr_translator:reset, fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_0_to_1_in_translator:reset, fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:reset, fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_0_to_2:wrreset_n, fifo_0_to_2_in_csr_translator:reset, fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_0_to_2_in_translator:reset, fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:reset, fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_1_to_0:rdreset_n, fifo_1_to_0_out_csr_translator:reset, fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:reset, fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_1_to_0_out_translator:reset, fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:reset, fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_2_to_0:rdreset_n, fifo_2_to_0_out_csr_translator:reset, fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:reset, fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_2_to_0_out_translator:reset, fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:reset, fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_003:reset, id_router_004:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_023:reset, id_router_024:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory_0:reset, onchip_memory_0_s1_translator:reset, onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, performance_counter_0:reset_n, performance_counter_0_control_slave_translator:reset, performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:reset, performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, timer_0_0:reset_n, timer_0_0_s1_translator:reset, timer_0_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0_1:reset_n, timer_0_1_s1_translator:reset, timer_0_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         rst_controller_reset_out_reset_req;                                                                       // rst_controller:reset_req -> onchip_memory_0:reset_req
	wire         cpu_0_jtag_debug_module_reset_reset;                                                                      // cpu_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller_002:reset_in0]
	wire         rst_controller_001_reset_out_reset;                                                                       // rst_controller_001:reset_out -> [addr_router_002:reset, addr_router_003:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_mux_026:reset, cmd_xbar_mux_027:reset, cpu_1:reset_n, cpu_1_data_master_translator:reset, cpu_1_data_master_translator_avalon_universal_master_0_agent:reset, cpu_1_instruction_master_translator:reset, cpu_1_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_1_jtag_debug_module_translator:reset, cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_0_to_1:rdreset_n, fifo_0_to_1_out_csr_translator:reset, fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:reset, fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_0_to_1_out_translator:reset, fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:reset, fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_1_to_0:wrreset_n, fifo_1_to_0_in_csr_translator:reset, fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_1_to_0_in_translator:reset, fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:reset, fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_1_to_2:wrreset_n, fifo_1_to_2_in_csr_translator:reset, fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_1_to_2_in_translator:reset, fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:reset, fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_2_to_1:rdreset_n, fifo_2_to_1_out_csr_translator:reset, fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:reset, fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_2_to_1_out_translator:reset, fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:reset, fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_026:reset, id_router_027:reset, id_router_028:reset, id_router_029:reset, id_router_030:reset, id_router_031:reset, id_router_032:reset, id_router_033:reset, id_router_034:reset, id_router_035:reset, id_router_036:reset, id_router_037:reset, id_router_038:reset, id_router_039:reset, irq_mapper_001:reset, jtag_uart_1:rst_n, jtag_uart_1_avalon_jtag_slave_translator:reset, jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory_1:reset, onchip_memory_1_s1_translator:reset, onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, performance_counter_1:reset_n, performance_counter_1_control_slave_translator:reset, performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:reset, performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_026:reset, rsp_xbar_demux_027:reset, rsp_xbar_demux_028:reset, rsp_xbar_demux_029:reset, rsp_xbar_demux_030:reset, rsp_xbar_demux_031:reset, rsp_xbar_demux_032:reset, rsp_xbar_demux_033:reset, rsp_xbar_demux_034:reset, rsp_xbar_demux_035:reset, rsp_xbar_demux_036:reset, rsp_xbar_demux_037:reset, rsp_xbar_demux_038:reset, rsp_xbar_demux_039:reset, rsp_xbar_mux_002:reset, rsp_xbar_mux_003:reset, timer_1_0:reset_n, timer_1_0_s1_translator:reset, timer_1_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_1_1:reset_n, timer_1_1_s1_translator:reset, timer_1_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         rst_controller_001_reset_out_reset_req;                                                                   // rst_controller_001:reset_req -> onchip_memory_1:reset_req
	wire         cpu_1_jtag_debug_module_reset_reset;                                                                      // cpu_1:jtag_debug_module_resetrequest -> [rst_controller_001:reset_in0, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                                                                       // rst_controller_002:reset_out -> [cmd_xbar_mux_002:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, cmd_xbar_mux_007:reset, cmd_xbar_mux_008:reset, cmd_xbar_mux_009:reset, cmd_xbar_mux_010:reset, cmd_xbar_mux_019:reset, cmd_xbar_mux_020:reset, cmd_xbar_mux_021:reset, cmd_xbar_mux_022:reset, cmd_xbar_mux_025:reset, green_leds:reset_n, green_leds_s1_translator:reset, green_leds_s1_translator_avalon_universal_slave_0_agent:reset, green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_002:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, id_router_025:reset, mutex_0:reset_n, mutex_0_s1_translator:reset, mutex_0_s1_translator_avalon_universal_slave_0_agent:reset, mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, mutex_1:reset_n, mutex_1_s1_translator:reset, mutex_1_s1_translator_avalon_universal_slave_0_agent:reset, mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, mutex_2:reset_n, mutex_2_s1_translator:reset, mutex_2_s1_translator_avalon_universal_slave_0_agent:reset, mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, mutex_3:reset_n, mutex_3_s1_translator:reset, mutex_3_s1_translator_avalon_universal_slave_0_agent:reset, mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, mutex_4:reset_n, mutex_4_s1_translator:reset, mutex_4_s1_translator_avalon_universal_slave_0_agent:reset, mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, mutex_5:reset_n, mutex_5_s1_translator:reset, mutex_5_s1_translator_avalon_universal_slave_0_agent:reset, mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_shared:reset, onchip_shared_s1_translator:reset, onchip_shared_s1_translator_avalon_universal_slave_0_agent:reset, onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, red_leds:reset_n, red_leds_s1_translator:reset, red_leds_s1_translator_avalon_universal_slave_0_agent:reset, red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_025:reset, switches:reset_n, switches_s1_translator:reset, switches_s1_translator_avalon_universal_slave_0_agent:reset, switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_shared_0:reset_n, timer_shared_0_s1_translator:reset, timer_shared_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_shared_1:reset_n, timer_shared_1_s1_translator:reset, timer_shared_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         rst_controller_002_reset_out_reset_req;                                                                   // rst_controller_002:reset_req -> onchip_shared:reset_req
	wire         cpu_2_jtag_debug_module_reset_reset;                                                                      // cpu_2:jtag_debug_module_resetrequest -> [rst_controller_002:reset_in2, rst_controller_003:reset_in0]
	wire         rst_controller_003_reset_out_reset;                                                                       // rst_controller_003:reset_out -> [addr_router_004:reset, addr_router_005:reset, cmd_xbar_demux_004:reset, cmd_xbar_demux_005:reset, cmd_xbar_mux_040:reset, cmd_xbar_mux_041:reset, cpu_2:reset_n, cpu_2_data_master_translator:reset, cpu_2_data_master_translator_avalon_universal_master_0_agent:reset, cpu_2_instruction_master_translator:reset, cpu_2_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_2_jtag_debug_module_translator:reset, cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_0_to_2:rdreset_n, fifo_0_to_2_out_csr_translator:reset, fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:reset, fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_0_to_2_out_translator:reset, fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:reset, fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_1_to_2:rdreset_n, fifo_1_to_2_out_csr_translator:reset, fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:reset, fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_1_to_2_out_translator:reset, fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:reset, fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_2_to_0:wrreset_n, fifo_2_to_0_in_csr_translator:reset, fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_2_to_0_in_translator:reset, fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:reset, fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_2_to_1:wrreset_n, fifo_2_to_1_in_csr_translator:reset, fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_2_to_1_in_translator:reset, fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:reset, fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_040:reset, id_router_041:reset, id_router_042:reset, id_router_043:reset, id_router_044:reset, id_router_045:reset, id_router_046:reset, id_router_047:reset, id_router_048:reset, id_router_049:reset, id_router_050:reset, id_router_051:reset, id_router_052:reset, id_router_053:reset, irq_mapper_002:reset, jtag_uart_2:rst_n, jtag_uart_2_avalon_jtag_slave_translator:reset, jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory_2:reset, onchip_memory_2_s1_translator:reset, onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, performance_counter_2:reset_n, performance_counter_2_control_slave_translator:reset, performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:reset, performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_040:reset, rsp_xbar_demux_041:reset, rsp_xbar_demux_042:reset, rsp_xbar_demux_043:reset, rsp_xbar_demux_044:reset, rsp_xbar_demux_045:reset, rsp_xbar_demux_046:reset, rsp_xbar_demux_047:reset, rsp_xbar_demux_048:reset, rsp_xbar_demux_049:reset, rsp_xbar_demux_050:reset, rsp_xbar_demux_051:reset, rsp_xbar_demux_052:reset, rsp_xbar_demux_053:reset, rsp_xbar_mux_004:reset, rsp_xbar_mux_005:reset, timer_2_0:reset_n, timer_2_0_s1_translator:reset, timer_2_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_2_1:reset_n, timer_2_1_s1_translator:reset, timer_2_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         rst_controller_003_reset_out_reset_req;                                                                   // rst_controller_003:reset_req -> onchip_memory_2:reset_req
	wire         cmd_xbar_demux_src0_endofpacket;                                                                          // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                                // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                        // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_src0_data;                                                                                 // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire  [53:0] cmd_xbar_demux_src0_channel;                                                                              // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                                // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                          // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                                // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                        // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_src1_data;                                                                                 // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire  [53:0] cmd_xbar_demux_src1_channel;                                                                              // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                                // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                          // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                                // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                        // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_src2_data;                                                                                 // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire  [53:0] cmd_xbar_demux_src2_channel;                                                                              // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                                // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                      // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                            // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                                    // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src0_data;                                                                             // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire  [53:0] cmd_xbar_demux_001_src0_channel;                                                                          // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                            // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                      // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                            // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                                    // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src1_data;                                                                             // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire  [53:0] cmd_xbar_demux_001_src1_channel;                                                                          // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                            // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                      // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                            // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                                    // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src2_data;                                                                             // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire  [53:0] cmd_xbar_demux_001_src2_channel;                                                                          // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                            // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                      // cmd_xbar_demux_001:src3_endofpacket -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                            // cmd_xbar_demux_001:src3_valid -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                                    // cmd_xbar_demux_001:src3_startofpacket -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src3_data;                                                                             // cmd_xbar_demux_001:src3_data -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_001_src3_channel;                                                                          // cmd_xbar_demux_001:src3_channel -> timer_0_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                      // cmd_xbar_demux_001:src4_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                            // cmd_xbar_demux_001:src4_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                                    // cmd_xbar_demux_001:src4_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src4_data;                                                                             // cmd_xbar_demux_001:src4_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_001_src4_channel;                                                                          // cmd_xbar_demux_001:src4_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                      // cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                            // cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                                    // cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src5_data;                                                                             // cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink0_data
	wire  [53:0] cmd_xbar_demux_001_src5_channel;                                                                          // cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire         cmd_xbar_demux_001_src5_ready;                                                                            // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux_001:src5_ready
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                      // cmd_xbar_demux_001:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                            // cmd_xbar_demux_001:src6_valid -> cmd_xbar_mux_006:sink0_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                                    // cmd_xbar_demux_001:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src6_data;                                                                             // cmd_xbar_demux_001:src6_data -> cmd_xbar_mux_006:sink0_data
	wire  [53:0] cmd_xbar_demux_001_src6_channel;                                                                          // cmd_xbar_demux_001:src6_channel -> cmd_xbar_mux_006:sink0_channel
	wire         cmd_xbar_demux_001_src6_ready;                                                                            // cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux_001:src6_ready
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                      // cmd_xbar_demux_001:src7_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                            // cmd_xbar_demux_001:src7_valid -> cmd_xbar_mux_007:sink0_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                                    // cmd_xbar_demux_001:src7_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src7_data;                                                                             // cmd_xbar_demux_001:src7_data -> cmd_xbar_mux_007:sink0_data
	wire  [53:0] cmd_xbar_demux_001_src7_channel;                                                                          // cmd_xbar_demux_001:src7_channel -> cmd_xbar_mux_007:sink0_channel
	wire         cmd_xbar_demux_001_src7_ready;                                                                            // cmd_xbar_mux_007:sink0_ready -> cmd_xbar_demux_001:src7_ready
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                                      // cmd_xbar_demux_001:src8_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                            // cmd_xbar_demux_001:src8_valid -> cmd_xbar_mux_008:sink0_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                                    // cmd_xbar_demux_001:src8_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src8_data;                                                                             // cmd_xbar_demux_001:src8_data -> cmd_xbar_mux_008:sink0_data
	wire  [53:0] cmd_xbar_demux_001_src8_channel;                                                                          // cmd_xbar_demux_001:src8_channel -> cmd_xbar_mux_008:sink0_channel
	wire         cmd_xbar_demux_001_src8_ready;                                                                            // cmd_xbar_mux_008:sink0_ready -> cmd_xbar_demux_001:src8_ready
	wire         cmd_xbar_demux_001_src9_endofpacket;                                                                      // cmd_xbar_demux_001:src9_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	wire         cmd_xbar_demux_001_src9_valid;                                                                            // cmd_xbar_demux_001:src9_valid -> cmd_xbar_mux_009:sink0_valid
	wire         cmd_xbar_demux_001_src9_startofpacket;                                                                    // cmd_xbar_demux_001:src9_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src9_data;                                                                             // cmd_xbar_demux_001:src9_data -> cmd_xbar_mux_009:sink0_data
	wire  [53:0] cmd_xbar_demux_001_src9_channel;                                                                          // cmd_xbar_demux_001:src9_channel -> cmd_xbar_mux_009:sink0_channel
	wire         cmd_xbar_demux_001_src9_ready;                                                                            // cmd_xbar_mux_009:sink0_ready -> cmd_xbar_demux_001:src9_ready
	wire         cmd_xbar_demux_001_src10_endofpacket;                                                                     // cmd_xbar_demux_001:src10_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	wire         cmd_xbar_demux_001_src10_valid;                                                                           // cmd_xbar_demux_001:src10_valid -> cmd_xbar_mux_010:sink0_valid
	wire         cmd_xbar_demux_001_src10_startofpacket;                                                                   // cmd_xbar_demux_001:src10_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src10_data;                                                                            // cmd_xbar_demux_001:src10_data -> cmd_xbar_mux_010:sink0_data
	wire  [53:0] cmd_xbar_demux_001_src10_channel;                                                                         // cmd_xbar_demux_001:src10_channel -> cmd_xbar_mux_010:sink0_channel
	wire         cmd_xbar_demux_001_src10_ready;                                                                           // cmd_xbar_mux_010:sink0_ready -> cmd_xbar_demux_001:src10_ready
	wire         cmd_xbar_demux_001_src11_endofpacket;                                                                     // cmd_xbar_demux_001:src11_endofpacket -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src11_valid;                                                                           // cmd_xbar_demux_001:src11_valid -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src11_startofpacket;                                                                   // cmd_xbar_demux_001:src11_startofpacket -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src11_data;                                                                            // cmd_xbar_demux_001:src11_data -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_001_src11_channel;                                                                         // cmd_xbar_demux_001:src11_channel -> fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src12_endofpacket;                                                                     // cmd_xbar_demux_001:src12_endofpacket -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src12_valid;                                                                           // cmd_xbar_demux_001:src12_valid -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src12_startofpacket;                                                                   // cmd_xbar_demux_001:src12_startofpacket -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src12_data;                                                                            // cmd_xbar_demux_001:src12_data -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_001_src12_channel;                                                                         // cmd_xbar_demux_001:src12_channel -> fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src13_endofpacket;                                                                     // cmd_xbar_demux_001:src13_endofpacket -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src13_valid;                                                                           // cmd_xbar_demux_001:src13_valid -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src13_startofpacket;                                                                   // cmd_xbar_demux_001:src13_startofpacket -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src13_data;                                                                            // cmd_xbar_demux_001:src13_data -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_001_src13_channel;                                                                         // cmd_xbar_demux_001:src13_channel -> fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src14_endofpacket;                                                                     // cmd_xbar_demux_001:src14_endofpacket -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src14_valid;                                                                           // cmd_xbar_demux_001:src14_valid -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src14_startofpacket;                                                                   // cmd_xbar_demux_001:src14_startofpacket -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src14_data;                                                                            // cmd_xbar_demux_001:src14_data -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_001_src14_channel;                                                                         // cmd_xbar_demux_001:src14_channel -> fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src15_endofpacket;                                                                     // cmd_xbar_demux_001:src15_endofpacket -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src15_valid;                                                                           // cmd_xbar_demux_001:src15_valid -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src15_startofpacket;                                                                   // cmd_xbar_demux_001:src15_startofpacket -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src15_data;                                                                            // cmd_xbar_demux_001:src15_data -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_001_src15_channel;                                                                         // cmd_xbar_demux_001:src15_channel -> fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src16_endofpacket;                                                                     // cmd_xbar_demux_001:src16_endofpacket -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src16_valid;                                                                           // cmd_xbar_demux_001:src16_valid -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src16_startofpacket;                                                                   // cmd_xbar_demux_001:src16_startofpacket -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src16_data;                                                                            // cmd_xbar_demux_001:src16_data -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_001_src16_channel;                                                                         // cmd_xbar_demux_001:src16_channel -> fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src17_endofpacket;                                                                     // cmd_xbar_demux_001:src17_endofpacket -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src17_valid;                                                                           // cmd_xbar_demux_001:src17_valid -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src17_startofpacket;                                                                   // cmd_xbar_demux_001:src17_startofpacket -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src17_data;                                                                            // cmd_xbar_demux_001:src17_data -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_001_src17_channel;                                                                         // cmd_xbar_demux_001:src17_channel -> fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src18_endofpacket;                                                                     // cmd_xbar_demux_001:src18_endofpacket -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src18_valid;                                                                           // cmd_xbar_demux_001:src18_valid -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src18_startofpacket;                                                                   // cmd_xbar_demux_001:src18_startofpacket -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src18_data;                                                                            // cmd_xbar_demux_001:src18_data -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_001_src18_channel;                                                                         // cmd_xbar_demux_001:src18_channel -> fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src19_endofpacket;                                                                     // cmd_xbar_demux_001:src19_endofpacket -> cmd_xbar_mux_019:sink0_endofpacket
	wire         cmd_xbar_demux_001_src19_valid;                                                                           // cmd_xbar_demux_001:src19_valid -> cmd_xbar_mux_019:sink0_valid
	wire         cmd_xbar_demux_001_src19_startofpacket;                                                                   // cmd_xbar_demux_001:src19_startofpacket -> cmd_xbar_mux_019:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src19_data;                                                                            // cmd_xbar_demux_001:src19_data -> cmd_xbar_mux_019:sink0_data
	wire  [53:0] cmd_xbar_demux_001_src19_channel;                                                                         // cmd_xbar_demux_001:src19_channel -> cmd_xbar_mux_019:sink0_channel
	wire         cmd_xbar_demux_001_src19_ready;                                                                           // cmd_xbar_mux_019:sink0_ready -> cmd_xbar_demux_001:src19_ready
	wire         cmd_xbar_demux_001_src20_endofpacket;                                                                     // cmd_xbar_demux_001:src20_endofpacket -> cmd_xbar_mux_020:sink0_endofpacket
	wire         cmd_xbar_demux_001_src20_valid;                                                                           // cmd_xbar_demux_001:src20_valid -> cmd_xbar_mux_020:sink0_valid
	wire         cmd_xbar_demux_001_src20_startofpacket;                                                                   // cmd_xbar_demux_001:src20_startofpacket -> cmd_xbar_mux_020:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src20_data;                                                                            // cmd_xbar_demux_001:src20_data -> cmd_xbar_mux_020:sink0_data
	wire  [53:0] cmd_xbar_demux_001_src20_channel;                                                                         // cmd_xbar_demux_001:src20_channel -> cmd_xbar_mux_020:sink0_channel
	wire         cmd_xbar_demux_001_src20_ready;                                                                           // cmd_xbar_mux_020:sink0_ready -> cmd_xbar_demux_001:src20_ready
	wire         cmd_xbar_demux_001_src21_endofpacket;                                                                     // cmd_xbar_demux_001:src21_endofpacket -> cmd_xbar_mux_021:sink0_endofpacket
	wire         cmd_xbar_demux_001_src21_valid;                                                                           // cmd_xbar_demux_001:src21_valid -> cmd_xbar_mux_021:sink0_valid
	wire         cmd_xbar_demux_001_src21_startofpacket;                                                                   // cmd_xbar_demux_001:src21_startofpacket -> cmd_xbar_mux_021:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src21_data;                                                                            // cmd_xbar_demux_001:src21_data -> cmd_xbar_mux_021:sink0_data
	wire  [53:0] cmd_xbar_demux_001_src21_channel;                                                                         // cmd_xbar_demux_001:src21_channel -> cmd_xbar_mux_021:sink0_channel
	wire         cmd_xbar_demux_001_src21_ready;                                                                           // cmd_xbar_mux_021:sink0_ready -> cmd_xbar_demux_001:src21_ready
	wire         cmd_xbar_demux_001_src22_endofpacket;                                                                     // cmd_xbar_demux_001:src22_endofpacket -> cmd_xbar_mux_022:sink0_endofpacket
	wire         cmd_xbar_demux_001_src22_valid;                                                                           // cmd_xbar_demux_001:src22_valid -> cmd_xbar_mux_022:sink0_valid
	wire         cmd_xbar_demux_001_src22_startofpacket;                                                                   // cmd_xbar_demux_001:src22_startofpacket -> cmd_xbar_mux_022:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src22_data;                                                                            // cmd_xbar_demux_001:src22_data -> cmd_xbar_mux_022:sink0_data
	wire  [53:0] cmd_xbar_demux_001_src22_channel;                                                                         // cmd_xbar_demux_001:src22_channel -> cmd_xbar_mux_022:sink0_channel
	wire         cmd_xbar_demux_001_src22_ready;                                                                           // cmd_xbar_mux_022:sink0_ready -> cmd_xbar_demux_001:src22_ready
	wire         cmd_xbar_demux_001_src23_endofpacket;                                                                     // cmd_xbar_demux_001:src23_endofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src23_valid;                                                                           // cmd_xbar_demux_001:src23_valid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src23_startofpacket;                                                                   // cmd_xbar_demux_001:src23_startofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src23_data;                                                                            // cmd_xbar_demux_001:src23_data -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_001_src23_channel;                                                                         // cmd_xbar_demux_001:src23_channel -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src24_endofpacket;                                                                     // cmd_xbar_demux_001:src24_endofpacket -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src24_valid;                                                                           // cmd_xbar_demux_001:src24_valid -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src24_startofpacket;                                                                   // cmd_xbar_demux_001:src24_startofpacket -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src24_data;                                                                            // cmd_xbar_demux_001:src24_data -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_001_src24_channel;                                                                         // cmd_xbar_demux_001:src24_channel -> timer_0_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src25_endofpacket;                                                                     // cmd_xbar_demux_001:src25_endofpacket -> cmd_xbar_mux_025:sink0_endofpacket
	wire         cmd_xbar_demux_001_src25_valid;                                                                           // cmd_xbar_demux_001:src25_valid -> cmd_xbar_mux_025:sink0_valid
	wire         cmd_xbar_demux_001_src25_startofpacket;                                                                   // cmd_xbar_demux_001:src25_startofpacket -> cmd_xbar_mux_025:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_001_src25_data;                                                                            // cmd_xbar_demux_001:src25_data -> cmd_xbar_mux_025:sink0_data
	wire  [53:0] cmd_xbar_demux_001_src25_channel;                                                                         // cmd_xbar_demux_001:src25_channel -> cmd_xbar_mux_025:sink0_channel
	wire         cmd_xbar_demux_001_src25_ready;                                                                           // cmd_xbar_mux_025:sink0_ready -> cmd_xbar_demux_001:src25_ready
	wire         cmd_xbar_demux_002_src0_endofpacket;                                                                      // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_002:sink2_endofpacket
	wire         cmd_xbar_demux_002_src0_valid;                                                                            // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_002:sink2_valid
	wire         cmd_xbar_demux_002_src0_startofpacket;                                                                    // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_002:sink2_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src0_data;                                                                             // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_002:sink2_data
	wire  [53:0] cmd_xbar_demux_002_src0_channel;                                                                          // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_002:sink2_channel
	wire         cmd_xbar_demux_002_src0_ready;                                                                            // cmd_xbar_mux_002:sink2_ready -> cmd_xbar_demux_002:src0_ready
	wire         cmd_xbar_demux_002_src1_endofpacket;                                                                      // cmd_xbar_demux_002:src1_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire         cmd_xbar_demux_002_src1_valid;                                                                            // cmd_xbar_demux_002:src1_valid -> cmd_xbar_mux_005:sink1_valid
	wire         cmd_xbar_demux_002_src1_startofpacket;                                                                    // cmd_xbar_demux_002:src1_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src1_data;                                                                             // cmd_xbar_demux_002:src1_data -> cmd_xbar_mux_005:sink1_data
	wire  [53:0] cmd_xbar_demux_002_src1_channel;                                                                          // cmd_xbar_demux_002:src1_channel -> cmd_xbar_mux_005:sink1_channel
	wire         cmd_xbar_demux_002_src1_ready;                                                                            // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_002:src1_ready
	wire         cmd_xbar_demux_002_src2_endofpacket;                                                                      // cmd_xbar_demux_002:src2_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	wire         cmd_xbar_demux_002_src2_valid;                                                                            // cmd_xbar_demux_002:src2_valid -> cmd_xbar_mux_006:sink1_valid
	wire         cmd_xbar_demux_002_src2_startofpacket;                                                                    // cmd_xbar_demux_002:src2_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src2_data;                                                                             // cmd_xbar_demux_002:src2_data -> cmd_xbar_mux_006:sink1_data
	wire  [53:0] cmd_xbar_demux_002_src2_channel;                                                                          // cmd_xbar_demux_002:src2_channel -> cmd_xbar_mux_006:sink1_channel
	wire         cmd_xbar_demux_002_src2_ready;                                                                            // cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_002:src2_ready
	wire         cmd_xbar_demux_002_src3_endofpacket;                                                                      // cmd_xbar_demux_002:src3_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	wire         cmd_xbar_demux_002_src3_valid;                                                                            // cmd_xbar_demux_002:src3_valid -> cmd_xbar_mux_007:sink1_valid
	wire         cmd_xbar_demux_002_src3_startofpacket;                                                                    // cmd_xbar_demux_002:src3_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src3_data;                                                                             // cmd_xbar_demux_002:src3_data -> cmd_xbar_mux_007:sink1_data
	wire  [53:0] cmd_xbar_demux_002_src3_channel;                                                                          // cmd_xbar_demux_002:src3_channel -> cmd_xbar_mux_007:sink1_channel
	wire         cmd_xbar_demux_002_src3_ready;                                                                            // cmd_xbar_mux_007:sink1_ready -> cmd_xbar_demux_002:src3_ready
	wire         cmd_xbar_demux_002_src4_endofpacket;                                                                      // cmd_xbar_demux_002:src4_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	wire         cmd_xbar_demux_002_src4_valid;                                                                            // cmd_xbar_demux_002:src4_valid -> cmd_xbar_mux_008:sink1_valid
	wire         cmd_xbar_demux_002_src4_startofpacket;                                                                    // cmd_xbar_demux_002:src4_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src4_data;                                                                             // cmd_xbar_demux_002:src4_data -> cmd_xbar_mux_008:sink1_data
	wire  [53:0] cmd_xbar_demux_002_src4_channel;                                                                          // cmd_xbar_demux_002:src4_channel -> cmd_xbar_mux_008:sink1_channel
	wire         cmd_xbar_demux_002_src4_ready;                                                                            // cmd_xbar_mux_008:sink1_ready -> cmd_xbar_demux_002:src4_ready
	wire         cmd_xbar_demux_002_src5_endofpacket;                                                                      // cmd_xbar_demux_002:src5_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	wire         cmd_xbar_demux_002_src5_valid;                                                                            // cmd_xbar_demux_002:src5_valid -> cmd_xbar_mux_009:sink1_valid
	wire         cmd_xbar_demux_002_src5_startofpacket;                                                                    // cmd_xbar_demux_002:src5_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src5_data;                                                                             // cmd_xbar_demux_002:src5_data -> cmd_xbar_mux_009:sink1_data
	wire  [53:0] cmd_xbar_demux_002_src5_channel;                                                                          // cmd_xbar_demux_002:src5_channel -> cmd_xbar_mux_009:sink1_channel
	wire         cmd_xbar_demux_002_src5_ready;                                                                            // cmd_xbar_mux_009:sink1_ready -> cmd_xbar_demux_002:src5_ready
	wire         cmd_xbar_demux_002_src6_endofpacket;                                                                      // cmd_xbar_demux_002:src6_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	wire         cmd_xbar_demux_002_src6_valid;                                                                            // cmd_xbar_demux_002:src6_valid -> cmd_xbar_mux_010:sink1_valid
	wire         cmd_xbar_demux_002_src6_startofpacket;                                                                    // cmd_xbar_demux_002:src6_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src6_data;                                                                             // cmd_xbar_demux_002:src6_data -> cmd_xbar_mux_010:sink1_data
	wire  [53:0] cmd_xbar_demux_002_src6_channel;                                                                          // cmd_xbar_demux_002:src6_channel -> cmd_xbar_mux_010:sink1_channel
	wire         cmd_xbar_demux_002_src6_ready;                                                                            // cmd_xbar_mux_010:sink1_ready -> cmd_xbar_demux_002:src6_ready
	wire         cmd_xbar_demux_002_src7_endofpacket;                                                                      // cmd_xbar_demux_002:src7_endofpacket -> cmd_xbar_mux_019:sink1_endofpacket
	wire         cmd_xbar_demux_002_src7_valid;                                                                            // cmd_xbar_demux_002:src7_valid -> cmd_xbar_mux_019:sink1_valid
	wire         cmd_xbar_demux_002_src7_startofpacket;                                                                    // cmd_xbar_demux_002:src7_startofpacket -> cmd_xbar_mux_019:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src7_data;                                                                             // cmd_xbar_demux_002:src7_data -> cmd_xbar_mux_019:sink1_data
	wire  [53:0] cmd_xbar_demux_002_src7_channel;                                                                          // cmd_xbar_demux_002:src7_channel -> cmd_xbar_mux_019:sink1_channel
	wire         cmd_xbar_demux_002_src7_ready;                                                                            // cmd_xbar_mux_019:sink1_ready -> cmd_xbar_demux_002:src7_ready
	wire         cmd_xbar_demux_002_src8_endofpacket;                                                                      // cmd_xbar_demux_002:src8_endofpacket -> cmd_xbar_mux_020:sink1_endofpacket
	wire         cmd_xbar_demux_002_src8_valid;                                                                            // cmd_xbar_demux_002:src8_valid -> cmd_xbar_mux_020:sink1_valid
	wire         cmd_xbar_demux_002_src8_startofpacket;                                                                    // cmd_xbar_demux_002:src8_startofpacket -> cmd_xbar_mux_020:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src8_data;                                                                             // cmd_xbar_demux_002:src8_data -> cmd_xbar_mux_020:sink1_data
	wire  [53:0] cmd_xbar_demux_002_src8_channel;                                                                          // cmd_xbar_demux_002:src8_channel -> cmd_xbar_mux_020:sink1_channel
	wire         cmd_xbar_demux_002_src8_ready;                                                                            // cmd_xbar_mux_020:sink1_ready -> cmd_xbar_demux_002:src8_ready
	wire         cmd_xbar_demux_002_src9_endofpacket;                                                                      // cmd_xbar_demux_002:src9_endofpacket -> cmd_xbar_mux_021:sink1_endofpacket
	wire         cmd_xbar_demux_002_src9_valid;                                                                            // cmd_xbar_demux_002:src9_valid -> cmd_xbar_mux_021:sink1_valid
	wire         cmd_xbar_demux_002_src9_startofpacket;                                                                    // cmd_xbar_demux_002:src9_startofpacket -> cmd_xbar_mux_021:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src9_data;                                                                             // cmd_xbar_demux_002:src9_data -> cmd_xbar_mux_021:sink1_data
	wire  [53:0] cmd_xbar_demux_002_src9_channel;                                                                          // cmd_xbar_demux_002:src9_channel -> cmd_xbar_mux_021:sink1_channel
	wire         cmd_xbar_demux_002_src9_ready;                                                                            // cmd_xbar_mux_021:sink1_ready -> cmd_xbar_demux_002:src9_ready
	wire         cmd_xbar_demux_002_src10_endofpacket;                                                                     // cmd_xbar_demux_002:src10_endofpacket -> cmd_xbar_mux_022:sink1_endofpacket
	wire         cmd_xbar_demux_002_src10_valid;                                                                           // cmd_xbar_demux_002:src10_valid -> cmd_xbar_mux_022:sink1_valid
	wire         cmd_xbar_demux_002_src10_startofpacket;                                                                   // cmd_xbar_demux_002:src10_startofpacket -> cmd_xbar_mux_022:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src10_data;                                                                            // cmd_xbar_demux_002:src10_data -> cmd_xbar_mux_022:sink1_data
	wire  [53:0] cmd_xbar_demux_002_src10_channel;                                                                         // cmd_xbar_demux_002:src10_channel -> cmd_xbar_mux_022:sink1_channel
	wire         cmd_xbar_demux_002_src10_ready;                                                                           // cmd_xbar_mux_022:sink1_ready -> cmd_xbar_demux_002:src10_ready
	wire         cmd_xbar_demux_002_src11_endofpacket;                                                                     // cmd_xbar_demux_002:src11_endofpacket -> cmd_xbar_mux_025:sink1_endofpacket
	wire         cmd_xbar_demux_002_src11_valid;                                                                           // cmd_xbar_demux_002:src11_valid -> cmd_xbar_mux_025:sink1_valid
	wire         cmd_xbar_demux_002_src11_startofpacket;                                                                   // cmd_xbar_demux_002:src11_startofpacket -> cmd_xbar_mux_025:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src11_data;                                                                            // cmd_xbar_demux_002:src11_data -> cmd_xbar_mux_025:sink1_data
	wire  [53:0] cmd_xbar_demux_002_src11_channel;                                                                         // cmd_xbar_demux_002:src11_channel -> cmd_xbar_mux_025:sink1_channel
	wire         cmd_xbar_demux_002_src11_ready;                                                                           // cmd_xbar_mux_025:sink1_ready -> cmd_xbar_demux_002:src11_ready
	wire         cmd_xbar_demux_002_src12_endofpacket;                                                                     // cmd_xbar_demux_002:src12_endofpacket -> cmd_xbar_mux_026:sink0_endofpacket
	wire         cmd_xbar_demux_002_src12_valid;                                                                           // cmd_xbar_demux_002:src12_valid -> cmd_xbar_mux_026:sink0_valid
	wire         cmd_xbar_demux_002_src12_startofpacket;                                                                   // cmd_xbar_demux_002:src12_startofpacket -> cmd_xbar_mux_026:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src12_data;                                                                            // cmd_xbar_demux_002:src12_data -> cmd_xbar_mux_026:sink0_data
	wire  [53:0] cmd_xbar_demux_002_src12_channel;                                                                         // cmd_xbar_demux_002:src12_channel -> cmd_xbar_mux_026:sink0_channel
	wire         cmd_xbar_demux_002_src12_ready;                                                                           // cmd_xbar_mux_026:sink0_ready -> cmd_xbar_demux_002:src12_ready
	wire         cmd_xbar_demux_002_src13_endofpacket;                                                                     // cmd_xbar_demux_002:src13_endofpacket -> cmd_xbar_mux_027:sink0_endofpacket
	wire         cmd_xbar_demux_002_src13_valid;                                                                           // cmd_xbar_demux_002:src13_valid -> cmd_xbar_mux_027:sink0_valid
	wire         cmd_xbar_demux_002_src13_startofpacket;                                                                   // cmd_xbar_demux_002:src13_startofpacket -> cmd_xbar_mux_027:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src13_data;                                                                            // cmd_xbar_demux_002:src13_data -> cmd_xbar_mux_027:sink0_data
	wire  [53:0] cmd_xbar_demux_002_src13_channel;                                                                         // cmd_xbar_demux_002:src13_channel -> cmd_xbar_mux_027:sink0_channel
	wire         cmd_xbar_demux_002_src13_ready;                                                                           // cmd_xbar_mux_027:sink0_ready -> cmd_xbar_demux_002:src13_ready
	wire         cmd_xbar_demux_002_src14_endofpacket;                                                                     // cmd_xbar_demux_002:src14_endofpacket -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src14_valid;                                                                           // cmd_xbar_demux_002:src14_valid -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src14_startofpacket;                                                                   // cmd_xbar_demux_002:src14_startofpacket -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src14_data;                                                                            // cmd_xbar_demux_002:src14_data -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_002_src14_channel;                                                                         // cmd_xbar_demux_002:src14_channel -> timer_1_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src15_endofpacket;                                                                     // cmd_xbar_demux_002:src15_endofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src15_valid;                                                                           // cmd_xbar_demux_002:src15_valid -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src15_startofpacket;                                                                   // cmd_xbar_demux_002:src15_startofpacket -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src15_data;                                                                            // cmd_xbar_demux_002:src15_data -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_002_src15_channel;                                                                         // cmd_xbar_demux_002:src15_channel -> jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src16_endofpacket;                                                                     // cmd_xbar_demux_002:src16_endofpacket -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src16_valid;                                                                           // cmd_xbar_demux_002:src16_valid -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src16_startofpacket;                                                                   // cmd_xbar_demux_002:src16_startofpacket -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src16_data;                                                                            // cmd_xbar_demux_002:src16_data -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_002_src16_channel;                                                                         // cmd_xbar_demux_002:src16_channel -> fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src17_endofpacket;                                                                     // cmd_xbar_demux_002:src17_endofpacket -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src17_valid;                                                                           // cmd_xbar_demux_002:src17_valid -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src17_startofpacket;                                                                   // cmd_xbar_demux_002:src17_startofpacket -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src17_data;                                                                            // cmd_xbar_demux_002:src17_data -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_002_src17_channel;                                                                         // cmd_xbar_demux_002:src17_channel -> fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src18_endofpacket;                                                                     // cmd_xbar_demux_002:src18_endofpacket -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src18_valid;                                                                           // cmd_xbar_demux_002:src18_valid -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src18_startofpacket;                                                                   // cmd_xbar_demux_002:src18_startofpacket -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src18_data;                                                                            // cmd_xbar_demux_002:src18_data -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_002_src18_channel;                                                                         // cmd_xbar_demux_002:src18_channel -> fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src19_endofpacket;                                                                     // cmd_xbar_demux_002:src19_endofpacket -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src19_valid;                                                                           // cmd_xbar_demux_002:src19_valid -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src19_startofpacket;                                                                   // cmd_xbar_demux_002:src19_startofpacket -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src19_data;                                                                            // cmd_xbar_demux_002:src19_data -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_002_src19_channel;                                                                         // cmd_xbar_demux_002:src19_channel -> fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src20_endofpacket;                                                                     // cmd_xbar_demux_002:src20_endofpacket -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src20_valid;                                                                           // cmd_xbar_demux_002:src20_valid -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src20_startofpacket;                                                                   // cmd_xbar_demux_002:src20_startofpacket -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src20_data;                                                                            // cmd_xbar_demux_002:src20_data -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_002_src20_channel;                                                                         // cmd_xbar_demux_002:src20_channel -> fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src21_endofpacket;                                                                     // cmd_xbar_demux_002:src21_endofpacket -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src21_valid;                                                                           // cmd_xbar_demux_002:src21_valid -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src21_startofpacket;                                                                   // cmd_xbar_demux_002:src21_startofpacket -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src21_data;                                                                            // cmd_xbar_demux_002:src21_data -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_002_src21_channel;                                                                         // cmd_xbar_demux_002:src21_channel -> fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src22_endofpacket;                                                                     // cmd_xbar_demux_002:src22_endofpacket -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src22_valid;                                                                           // cmd_xbar_demux_002:src22_valid -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src22_startofpacket;                                                                   // cmd_xbar_demux_002:src22_startofpacket -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src22_data;                                                                            // cmd_xbar_demux_002:src22_data -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_002_src22_channel;                                                                         // cmd_xbar_demux_002:src22_channel -> fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src23_endofpacket;                                                                     // cmd_xbar_demux_002:src23_endofpacket -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src23_valid;                                                                           // cmd_xbar_demux_002:src23_valid -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src23_startofpacket;                                                                   // cmd_xbar_demux_002:src23_startofpacket -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src23_data;                                                                            // cmd_xbar_demux_002:src23_data -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_002_src23_channel;                                                                         // cmd_xbar_demux_002:src23_channel -> fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src24_endofpacket;                                                                     // cmd_xbar_demux_002:src24_endofpacket -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src24_valid;                                                                           // cmd_xbar_demux_002:src24_valid -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src24_startofpacket;                                                                   // cmd_xbar_demux_002:src24_startofpacket -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src24_data;                                                                            // cmd_xbar_demux_002:src24_data -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_002_src24_channel;                                                                         // cmd_xbar_demux_002:src24_channel -> performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src25_endofpacket;                                                                     // cmd_xbar_demux_002:src25_endofpacket -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_002_src25_valid;                                                                           // cmd_xbar_demux_002:src25_valid -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_002_src25_startofpacket;                                                                   // cmd_xbar_demux_002:src25_startofpacket -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_002_src25_data;                                                                            // cmd_xbar_demux_002:src25_data -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_002_src25_channel;                                                                         // cmd_xbar_demux_002:src25_channel -> timer_1_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_003_src0_endofpacket;                                                                      // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_002:sink3_endofpacket
	wire         cmd_xbar_demux_003_src0_valid;                                                                            // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_002:sink3_valid
	wire         cmd_xbar_demux_003_src0_startofpacket;                                                                    // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_002:sink3_startofpacket
	wire  [96:0] cmd_xbar_demux_003_src0_data;                                                                             // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_002:sink3_data
	wire  [53:0] cmd_xbar_demux_003_src0_channel;                                                                          // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_002:sink3_channel
	wire         cmd_xbar_demux_003_src0_ready;                                                                            // cmd_xbar_mux_002:sink3_ready -> cmd_xbar_demux_003:src0_ready
	wire         cmd_xbar_demux_003_src1_endofpacket;                                                                      // cmd_xbar_demux_003:src1_endofpacket -> cmd_xbar_mux_026:sink1_endofpacket
	wire         cmd_xbar_demux_003_src1_valid;                                                                            // cmd_xbar_demux_003:src1_valid -> cmd_xbar_mux_026:sink1_valid
	wire         cmd_xbar_demux_003_src1_startofpacket;                                                                    // cmd_xbar_demux_003:src1_startofpacket -> cmd_xbar_mux_026:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_003_src1_data;                                                                             // cmd_xbar_demux_003:src1_data -> cmd_xbar_mux_026:sink1_data
	wire  [53:0] cmd_xbar_demux_003_src1_channel;                                                                          // cmd_xbar_demux_003:src1_channel -> cmd_xbar_mux_026:sink1_channel
	wire         cmd_xbar_demux_003_src1_ready;                                                                            // cmd_xbar_mux_026:sink1_ready -> cmd_xbar_demux_003:src1_ready
	wire         cmd_xbar_demux_003_src2_endofpacket;                                                                      // cmd_xbar_demux_003:src2_endofpacket -> cmd_xbar_mux_027:sink1_endofpacket
	wire         cmd_xbar_demux_003_src2_valid;                                                                            // cmd_xbar_demux_003:src2_valid -> cmd_xbar_mux_027:sink1_valid
	wire         cmd_xbar_demux_003_src2_startofpacket;                                                                    // cmd_xbar_demux_003:src2_startofpacket -> cmd_xbar_mux_027:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_003_src2_data;                                                                             // cmd_xbar_demux_003:src2_data -> cmd_xbar_mux_027:sink1_data
	wire  [53:0] cmd_xbar_demux_003_src2_channel;                                                                          // cmd_xbar_demux_003:src2_channel -> cmd_xbar_mux_027:sink1_channel
	wire         cmd_xbar_demux_003_src2_ready;                                                                            // cmd_xbar_mux_027:sink1_ready -> cmd_xbar_demux_003:src2_ready
	wire         cmd_xbar_demux_004_src0_endofpacket;                                                                      // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_002:sink4_endofpacket
	wire         cmd_xbar_demux_004_src0_valid;                                                                            // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_002:sink4_valid
	wire         cmd_xbar_demux_004_src0_startofpacket;                                                                    // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_002:sink4_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src0_data;                                                                             // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_002:sink4_data
	wire  [53:0] cmd_xbar_demux_004_src0_channel;                                                                          // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_002:sink4_channel
	wire         cmd_xbar_demux_004_src0_ready;                                                                            // cmd_xbar_mux_002:sink4_ready -> cmd_xbar_demux_004:src0_ready
	wire         cmd_xbar_demux_004_src1_endofpacket;                                                                      // cmd_xbar_demux_004:src1_endofpacket -> cmd_xbar_mux_005:sink2_endofpacket
	wire         cmd_xbar_demux_004_src1_valid;                                                                            // cmd_xbar_demux_004:src1_valid -> cmd_xbar_mux_005:sink2_valid
	wire         cmd_xbar_demux_004_src1_startofpacket;                                                                    // cmd_xbar_demux_004:src1_startofpacket -> cmd_xbar_mux_005:sink2_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src1_data;                                                                             // cmd_xbar_demux_004:src1_data -> cmd_xbar_mux_005:sink2_data
	wire  [53:0] cmd_xbar_demux_004_src1_channel;                                                                          // cmd_xbar_demux_004:src1_channel -> cmd_xbar_mux_005:sink2_channel
	wire         cmd_xbar_demux_004_src1_ready;                                                                            // cmd_xbar_mux_005:sink2_ready -> cmd_xbar_demux_004:src1_ready
	wire         cmd_xbar_demux_004_src2_endofpacket;                                                                      // cmd_xbar_demux_004:src2_endofpacket -> cmd_xbar_mux_006:sink2_endofpacket
	wire         cmd_xbar_demux_004_src2_valid;                                                                            // cmd_xbar_demux_004:src2_valid -> cmd_xbar_mux_006:sink2_valid
	wire         cmd_xbar_demux_004_src2_startofpacket;                                                                    // cmd_xbar_demux_004:src2_startofpacket -> cmd_xbar_mux_006:sink2_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src2_data;                                                                             // cmd_xbar_demux_004:src2_data -> cmd_xbar_mux_006:sink2_data
	wire  [53:0] cmd_xbar_demux_004_src2_channel;                                                                          // cmd_xbar_demux_004:src2_channel -> cmd_xbar_mux_006:sink2_channel
	wire         cmd_xbar_demux_004_src2_ready;                                                                            // cmd_xbar_mux_006:sink2_ready -> cmd_xbar_demux_004:src2_ready
	wire         cmd_xbar_demux_004_src3_endofpacket;                                                                      // cmd_xbar_demux_004:src3_endofpacket -> cmd_xbar_mux_007:sink2_endofpacket
	wire         cmd_xbar_demux_004_src3_valid;                                                                            // cmd_xbar_demux_004:src3_valid -> cmd_xbar_mux_007:sink2_valid
	wire         cmd_xbar_demux_004_src3_startofpacket;                                                                    // cmd_xbar_demux_004:src3_startofpacket -> cmd_xbar_mux_007:sink2_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src3_data;                                                                             // cmd_xbar_demux_004:src3_data -> cmd_xbar_mux_007:sink2_data
	wire  [53:0] cmd_xbar_demux_004_src3_channel;                                                                          // cmd_xbar_demux_004:src3_channel -> cmd_xbar_mux_007:sink2_channel
	wire         cmd_xbar_demux_004_src3_ready;                                                                            // cmd_xbar_mux_007:sink2_ready -> cmd_xbar_demux_004:src3_ready
	wire         cmd_xbar_demux_004_src4_endofpacket;                                                                      // cmd_xbar_demux_004:src4_endofpacket -> cmd_xbar_mux_008:sink2_endofpacket
	wire         cmd_xbar_demux_004_src4_valid;                                                                            // cmd_xbar_demux_004:src4_valid -> cmd_xbar_mux_008:sink2_valid
	wire         cmd_xbar_demux_004_src4_startofpacket;                                                                    // cmd_xbar_demux_004:src4_startofpacket -> cmd_xbar_mux_008:sink2_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src4_data;                                                                             // cmd_xbar_demux_004:src4_data -> cmd_xbar_mux_008:sink2_data
	wire  [53:0] cmd_xbar_demux_004_src4_channel;                                                                          // cmd_xbar_demux_004:src4_channel -> cmd_xbar_mux_008:sink2_channel
	wire         cmd_xbar_demux_004_src4_ready;                                                                            // cmd_xbar_mux_008:sink2_ready -> cmd_xbar_demux_004:src4_ready
	wire         cmd_xbar_demux_004_src5_endofpacket;                                                                      // cmd_xbar_demux_004:src5_endofpacket -> cmd_xbar_mux_009:sink2_endofpacket
	wire         cmd_xbar_demux_004_src5_valid;                                                                            // cmd_xbar_demux_004:src5_valid -> cmd_xbar_mux_009:sink2_valid
	wire         cmd_xbar_demux_004_src5_startofpacket;                                                                    // cmd_xbar_demux_004:src5_startofpacket -> cmd_xbar_mux_009:sink2_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src5_data;                                                                             // cmd_xbar_demux_004:src5_data -> cmd_xbar_mux_009:sink2_data
	wire  [53:0] cmd_xbar_demux_004_src5_channel;                                                                          // cmd_xbar_demux_004:src5_channel -> cmd_xbar_mux_009:sink2_channel
	wire         cmd_xbar_demux_004_src5_ready;                                                                            // cmd_xbar_mux_009:sink2_ready -> cmd_xbar_demux_004:src5_ready
	wire         cmd_xbar_demux_004_src6_endofpacket;                                                                      // cmd_xbar_demux_004:src6_endofpacket -> cmd_xbar_mux_010:sink2_endofpacket
	wire         cmd_xbar_demux_004_src6_valid;                                                                            // cmd_xbar_demux_004:src6_valid -> cmd_xbar_mux_010:sink2_valid
	wire         cmd_xbar_demux_004_src6_startofpacket;                                                                    // cmd_xbar_demux_004:src6_startofpacket -> cmd_xbar_mux_010:sink2_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src6_data;                                                                             // cmd_xbar_demux_004:src6_data -> cmd_xbar_mux_010:sink2_data
	wire  [53:0] cmd_xbar_demux_004_src6_channel;                                                                          // cmd_xbar_demux_004:src6_channel -> cmd_xbar_mux_010:sink2_channel
	wire         cmd_xbar_demux_004_src6_ready;                                                                            // cmd_xbar_mux_010:sink2_ready -> cmd_xbar_demux_004:src6_ready
	wire         cmd_xbar_demux_004_src7_endofpacket;                                                                      // cmd_xbar_demux_004:src7_endofpacket -> cmd_xbar_mux_019:sink2_endofpacket
	wire         cmd_xbar_demux_004_src7_valid;                                                                            // cmd_xbar_demux_004:src7_valid -> cmd_xbar_mux_019:sink2_valid
	wire         cmd_xbar_demux_004_src7_startofpacket;                                                                    // cmd_xbar_demux_004:src7_startofpacket -> cmd_xbar_mux_019:sink2_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src7_data;                                                                             // cmd_xbar_demux_004:src7_data -> cmd_xbar_mux_019:sink2_data
	wire  [53:0] cmd_xbar_demux_004_src7_channel;                                                                          // cmd_xbar_demux_004:src7_channel -> cmd_xbar_mux_019:sink2_channel
	wire         cmd_xbar_demux_004_src7_ready;                                                                            // cmd_xbar_mux_019:sink2_ready -> cmd_xbar_demux_004:src7_ready
	wire         cmd_xbar_demux_004_src8_endofpacket;                                                                      // cmd_xbar_demux_004:src8_endofpacket -> cmd_xbar_mux_020:sink2_endofpacket
	wire         cmd_xbar_demux_004_src8_valid;                                                                            // cmd_xbar_demux_004:src8_valid -> cmd_xbar_mux_020:sink2_valid
	wire         cmd_xbar_demux_004_src8_startofpacket;                                                                    // cmd_xbar_demux_004:src8_startofpacket -> cmd_xbar_mux_020:sink2_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src8_data;                                                                             // cmd_xbar_demux_004:src8_data -> cmd_xbar_mux_020:sink2_data
	wire  [53:0] cmd_xbar_demux_004_src8_channel;                                                                          // cmd_xbar_demux_004:src8_channel -> cmd_xbar_mux_020:sink2_channel
	wire         cmd_xbar_demux_004_src8_ready;                                                                            // cmd_xbar_mux_020:sink2_ready -> cmd_xbar_demux_004:src8_ready
	wire         cmd_xbar_demux_004_src9_endofpacket;                                                                      // cmd_xbar_demux_004:src9_endofpacket -> cmd_xbar_mux_021:sink2_endofpacket
	wire         cmd_xbar_demux_004_src9_valid;                                                                            // cmd_xbar_demux_004:src9_valid -> cmd_xbar_mux_021:sink2_valid
	wire         cmd_xbar_demux_004_src9_startofpacket;                                                                    // cmd_xbar_demux_004:src9_startofpacket -> cmd_xbar_mux_021:sink2_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src9_data;                                                                             // cmd_xbar_demux_004:src9_data -> cmd_xbar_mux_021:sink2_data
	wire  [53:0] cmd_xbar_demux_004_src9_channel;                                                                          // cmd_xbar_demux_004:src9_channel -> cmd_xbar_mux_021:sink2_channel
	wire         cmd_xbar_demux_004_src9_ready;                                                                            // cmd_xbar_mux_021:sink2_ready -> cmd_xbar_demux_004:src9_ready
	wire         cmd_xbar_demux_004_src10_endofpacket;                                                                     // cmd_xbar_demux_004:src10_endofpacket -> cmd_xbar_mux_022:sink2_endofpacket
	wire         cmd_xbar_demux_004_src10_valid;                                                                           // cmd_xbar_demux_004:src10_valid -> cmd_xbar_mux_022:sink2_valid
	wire         cmd_xbar_demux_004_src10_startofpacket;                                                                   // cmd_xbar_demux_004:src10_startofpacket -> cmd_xbar_mux_022:sink2_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src10_data;                                                                            // cmd_xbar_demux_004:src10_data -> cmd_xbar_mux_022:sink2_data
	wire  [53:0] cmd_xbar_demux_004_src10_channel;                                                                         // cmd_xbar_demux_004:src10_channel -> cmd_xbar_mux_022:sink2_channel
	wire         cmd_xbar_demux_004_src10_ready;                                                                           // cmd_xbar_mux_022:sink2_ready -> cmd_xbar_demux_004:src10_ready
	wire         cmd_xbar_demux_004_src11_endofpacket;                                                                     // cmd_xbar_demux_004:src11_endofpacket -> cmd_xbar_mux_025:sink2_endofpacket
	wire         cmd_xbar_demux_004_src11_valid;                                                                           // cmd_xbar_demux_004:src11_valid -> cmd_xbar_mux_025:sink2_valid
	wire         cmd_xbar_demux_004_src11_startofpacket;                                                                   // cmd_xbar_demux_004:src11_startofpacket -> cmd_xbar_mux_025:sink2_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src11_data;                                                                            // cmd_xbar_demux_004:src11_data -> cmd_xbar_mux_025:sink2_data
	wire  [53:0] cmd_xbar_demux_004_src11_channel;                                                                         // cmd_xbar_demux_004:src11_channel -> cmd_xbar_mux_025:sink2_channel
	wire         cmd_xbar_demux_004_src11_ready;                                                                           // cmd_xbar_mux_025:sink2_ready -> cmd_xbar_demux_004:src11_ready
	wire         cmd_xbar_demux_004_src12_endofpacket;                                                                     // cmd_xbar_demux_004:src12_endofpacket -> cmd_xbar_mux_040:sink0_endofpacket
	wire         cmd_xbar_demux_004_src12_valid;                                                                           // cmd_xbar_demux_004:src12_valid -> cmd_xbar_mux_040:sink0_valid
	wire         cmd_xbar_demux_004_src12_startofpacket;                                                                   // cmd_xbar_demux_004:src12_startofpacket -> cmd_xbar_mux_040:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src12_data;                                                                            // cmd_xbar_demux_004:src12_data -> cmd_xbar_mux_040:sink0_data
	wire  [53:0] cmd_xbar_demux_004_src12_channel;                                                                         // cmd_xbar_demux_004:src12_channel -> cmd_xbar_mux_040:sink0_channel
	wire         cmd_xbar_demux_004_src12_ready;                                                                           // cmd_xbar_mux_040:sink0_ready -> cmd_xbar_demux_004:src12_ready
	wire         cmd_xbar_demux_004_src13_endofpacket;                                                                     // cmd_xbar_demux_004:src13_endofpacket -> cmd_xbar_mux_041:sink0_endofpacket
	wire         cmd_xbar_demux_004_src13_valid;                                                                           // cmd_xbar_demux_004:src13_valid -> cmd_xbar_mux_041:sink0_valid
	wire         cmd_xbar_demux_004_src13_startofpacket;                                                                   // cmd_xbar_demux_004:src13_startofpacket -> cmd_xbar_mux_041:sink0_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src13_data;                                                                            // cmd_xbar_demux_004:src13_data -> cmd_xbar_mux_041:sink0_data
	wire  [53:0] cmd_xbar_demux_004_src13_channel;                                                                         // cmd_xbar_demux_004:src13_channel -> cmd_xbar_mux_041:sink0_channel
	wire         cmd_xbar_demux_004_src13_ready;                                                                           // cmd_xbar_mux_041:sink0_ready -> cmd_xbar_demux_004:src13_ready
	wire         cmd_xbar_demux_004_src14_endofpacket;                                                                     // cmd_xbar_demux_004:src14_endofpacket -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src14_valid;                                                                           // cmd_xbar_demux_004:src14_valid -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src14_startofpacket;                                                                   // cmd_xbar_demux_004:src14_startofpacket -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src14_data;                                                                            // cmd_xbar_demux_004:src14_data -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_004_src14_channel;                                                                         // cmd_xbar_demux_004:src14_channel -> timer_2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src15_endofpacket;                                                                     // cmd_xbar_demux_004:src15_endofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src15_valid;                                                                           // cmd_xbar_demux_004:src15_valid -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src15_startofpacket;                                                                   // cmd_xbar_demux_004:src15_startofpacket -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src15_data;                                                                            // cmd_xbar_demux_004:src15_data -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_004_src15_channel;                                                                         // cmd_xbar_demux_004:src15_channel -> jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src16_endofpacket;                                                                     // cmd_xbar_demux_004:src16_endofpacket -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src16_valid;                                                                           // cmd_xbar_demux_004:src16_valid -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src16_startofpacket;                                                                   // cmd_xbar_demux_004:src16_startofpacket -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src16_data;                                                                            // cmd_xbar_demux_004:src16_data -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_004_src16_channel;                                                                         // cmd_xbar_demux_004:src16_channel -> fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src17_endofpacket;                                                                     // cmd_xbar_demux_004:src17_endofpacket -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src17_valid;                                                                           // cmd_xbar_demux_004:src17_valid -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src17_startofpacket;                                                                   // cmd_xbar_demux_004:src17_startofpacket -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src17_data;                                                                            // cmd_xbar_demux_004:src17_data -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_004_src17_channel;                                                                         // cmd_xbar_demux_004:src17_channel -> fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src18_endofpacket;                                                                     // cmd_xbar_demux_004:src18_endofpacket -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src18_valid;                                                                           // cmd_xbar_demux_004:src18_valid -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src18_startofpacket;                                                                   // cmd_xbar_demux_004:src18_startofpacket -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src18_data;                                                                            // cmd_xbar_demux_004:src18_data -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_004_src18_channel;                                                                         // cmd_xbar_demux_004:src18_channel -> fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src19_endofpacket;                                                                     // cmd_xbar_demux_004:src19_endofpacket -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src19_valid;                                                                           // cmd_xbar_demux_004:src19_valid -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src19_startofpacket;                                                                   // cmd_xbar_demux_004:src19_startofpacket -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src19_data;                                                                            // cmd_xbar_demux_004:src19_data -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_004_src19_channel;                                                                         // cmd_xbar_demux_004:src19_channel -> fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src20_endofpacket;                                                                     // cmd_xbar_demux_004:src20_endofpacket -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src20_valid;                                                                           // cmd_xbar_demux_004:src20_valid -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src20_startofpacket;                                                                   // cmd_xbar_demux_004:src20_startofpacket -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src20_data;                                                                            // cmd_xbar_demux_004:src20_data -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_004_src20_channel;                                                                         // cmd_xbar_demux_004:src20_channel -> fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src21_endofpacket;                                                                     // cmd_xbar_demux_004:src21_endofpacket -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src21_valid;                                                                           // cmd_xbar_demux_004:src21_valid -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src21_startofpacket;                                                                   // cmd_xbar_demux_004:src21_startofpacket -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src21_data;                                                                            // cmd_xbar_demux_004:src21_data -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_004_src21_channel;                                                                         // cmd_xbar_demux_004:src21_channel -> fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src22_endofpacket;                                                                     // cmd_xbar_demux_004:src22_endofpacket -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src22_valid;                                                                           // cmd_xbar_demux_004:src22_valid -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src22_startofpacket;                                                                   // cmd_xbar_demux_004:src22_startofpacket -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src22_data;                                                                            // cmd_xbar_demux_004:src22_data -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_004_src22_channel;                                                                         // cmd_xbar_demux_004:src22_channel -> fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src23_endofpacket;                                                                     // cmd_xbar_demux_004:src23_endofpacket -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src23_valid;                                                                           // cmd_xbar_demux_004:src23_valid -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src23_startofpacket;                                                                   // cmd_xbar_demux_004:src23_startofpacket -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src23_data;                                                                            // cmd_xbar_demux_004:src23_data -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_004_src23_channel;                                                                         // cmd_xbar_demux_004:src23_channel -> fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src24_endofpacket;                                                                     // cmd_xbar_demux_004:src24_endofpacket -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src24_valid;                                                                           // cmd_xbar_demux_004:src24_valid -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src24_startofpacket;                                                                   // cmd_xbar_demux_004:src24_startofpacket -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src24_data;                                                                            // cmd_xbar_demux_004:src24_data -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_004_src24_channel;                                                                         // cmd_xbar_demux_004:src24_channel -> performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_004_src25_endofpacket;                                                                     // cmd_xbar_demux_004:src25_endofpacket -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_004_src25_valid;                                                                           // cmd_xbar_demux_004:src25_valid -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_004_src25_startofpacket;                                                                   // cmd_xbar_demux_004:src25_startofpacket -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_demux_004_src25_data;                                                                            // cmd_xbar_demux_004:src25_data -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_demux_004_src25_channel;                                                                         // cmd_xbar_demux_004:src25_channel -> timer_2_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_005_src0_endofpacket;                                                                      // cmd_xbar_demux_005:src0_endofpacket -> cmd_xbar_mux_002:sink5_endofpacket
	wire         cmd_xbar_demux_005_src0_valid;                                                                            // cmd_xbar_demux_005:src0_valid -> cmd_xbar_mux_002:sink5_valid
	wire         cmd_xbar_demux_005_src0_startofpacket;                                                                    // cmd_xbar_demux_005:src0_startofpacket -> cmd_xbar_mux_002:sink5_startofpacket
	wire  [96:0] cmd_xbar_demux_005_src0_data;                                                                             // cmd_xbar_demux_005:src0_data -> cmd_xbar_mux_002:sink5_data
	wire  [53:0] cmd_xbar_demux_005_src0_channel;                                                                          // cmd_xbar_demux_005:src0_channel -> cmd_xbar_mux_002:sink5_channel
	wire         cmd_xbar_demux_005_src0_ready;                                                                            // cmd_xbar_mux_002:sink5_ready -> cmd_xbar_demux_005:src0_ready
	wire         cmd_xbar_demux_005_src1_endofpacket;                                                                      // cmd_xbar_demux_005:src1_endofpacket -> cmd_xbar_mux_040:sink1_endofpacket
	wire         cmd_xbar_demux_005_src1_valid;                                                                            // cmd_xbar_demux_005:src1_valid -> cmd_xbar_mux_040:sink1_valid
	wire         cmd_xbar_demux_005_src1_startofpacket;                                                                    // cmd_xbar_demux_005:src1_startofpacket -> cmd_xbar_mux_040:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_005_src1_data;                                                                             // cmd_xbar_demux_005:src1_data -> cmd_xbar_mux_040:sink1_data
	wire  [53:0] cmd_xbar_demux_005_src1_channel;                                                                          // cmd_xbar_demux_005:src1_channel -> cmd_xbar_mux_040:sink1_channel
	wire         cmd_xbar_demux_005_src1_ready;                                                                            // cmd_xbar_mux_040:sink1_ready -> cmd_xbar_demux_005:src1_ready
	wire         cmd_xbar_demux_005_src2_endofpacket;                                                                      // cmd_xbar_demux_005:src2_endofpacket -> cmd_xbar_mux_041:sink1_endofpacket
	wire         cmd_xbar_demux_005_src2_valid;                                                                            // cmd_xbar_demux_005:src2_valid -> cmd_xbar_mux_041:sink1_valid
	wire         cmd_xbar_demux_005_src2_startofpacket;                                                                    // cmd_xbar_demux_005:src2_startofpacket -> cmd_xbar_mux_041:sink1_startofpacket
	wire  [96:0] cmd_xbar_demux_005_src2_data;                                                                             // cmd_xbar_demux_005:src2_data -> cmd_xbar_mux_041:sink1_data
	wire  [53:0] cmd_xbar_demux_005_src2_channel;                                                                          // cmd_xbar_demux_005:src2_channel -> cmd_xbar_mux_041:sink1_channel
	wire         cmd_xbar_demux_005_src2_ready;                                                                            // cmd_xbar_mux_041:sink1_ready -> cmd_xbar_demux_005:src2_ready
	wire         rsp_xbar_demux_src0_endofpacket;                                                                          // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                                // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                        // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [96:0] rsp_xbar_demux_src0_data;                                                                                 // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [53:0] rsp_xbar_demux_src0_channel;                                                                              // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                                // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                          // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                                // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                        // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [96:0] rsp_xbar_demux_src1_data;                                                                                 // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire  [53:0] rsp_xbar_demux_src1_channel;                                                                              // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                                // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                      // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                            // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                                    // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [96:0] rsp_xbar_demux_001_src0_data;                                                                             // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [53:0] rsp_xbar_demux_001_src0_channel;                                                                          // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                            // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                      // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                            // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                                    // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [96:0] rsp_xbar_demux_001_src1_data;                                                                             // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire  [53:0] rsp_xbar_demux_001_src1_channel;                                                                          // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                            // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                      // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                            // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                                    // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [96:0] rsp_xbar_demux_002_src0_data;                                                                             // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire  [53:0] rsp_xbar_demux_002_src0_channel;                                                                          // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                            // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                      // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                            // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                                    // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [96:0] rsp_xbar_demux_002_src1_data;                                                                             // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire  [53:0] rsp_xbar_demux_002_src1_channel;                                                                          // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                            // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_002_src2_endofpacket;                                                                      // rsp_xbar_demux_002:src2_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire         rsp_xbar_demux_002_src2_valid;                                                                            // rsp_xbar_demux_002:src2_valid -> rsp_xbar_mux_002:sink0_valid
	wire         rsp_xbar_demux_002_src2_startofpacket;                                                                    // rsp_xbar_demux_002:src2_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire  [96:0] rsp_xbar_demux_002_src2_data;                                                                             // rsp_xbar_demux_002:src2_data -> rsp_xbar_mux_002:sink0_data
	wire  [53:0] rsp_xbar_demux_002_src2_channel;                                                                          // rsp_xbar_demux_002:src2_channel -> rsp_xbar_mux_002:sink0_channel
	wire         rsp_xbar_demux_002_src2_ready;                                                                            // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux_002:src2_ready
	wire         rsp_xbar_demux_002_src3_endofpacket;                                                                      // rsp_xbar_demux_002:src3_endofpacket -> rsp_xbar_mux_003:sink0_endofpacket
	wire         rsp_xbar_demux_002_src3_valid;                                                                            // rsp_xbar_demux_002:src3_valid -> rsp_xbar_mux_003:sink0_valid
	wire         rsp_xbar_demux_002_src3_startofpacket;                                                                    // rsp_xbar_demux_002:src3_startofpacket -> rsp_xbar_mux_003:sink0_startofpacket
	wire  [96:0] rsp_xbar_demux_002_src3_data;                                                                             // rsp_xbar_demux_002:src3_data -> rsp_xbar_mux_003:sink0_data
	wire  [53:0] rsp_xbar_demux_002_src3_channel;                                                                          // rsp_xbar_demux_002:src3_channel -> rsp_xbar_mux_003:sink0_channel
	wire         rsp_xbar_demux_002_src3_ready;                                                                            // rsp_xbar_mux_003:sink0_ready -> rsp_xbar_demux_002:src3_ready
	wire         rsp_xbar_demux_002_src4_endofpacket;                                                                      // rsp_xbar_demux_002:src4_endofpacket -> rsp_xbar_mux_004:sink0_endofpacket
	wire         rsp_xbar_demux_002_src4_valid;                                                                            // rsp_xbar_demux_002:src4_valid -> rsp_xbar_mux_004:sink0_valid
	wire         rsp_xbar_demux_002_src4_startofpacket;                                                                    // rsp_xbar_demux_002:src4_startofpacket -> rsp_xbar_mux_004:sink0_startofpacket
	wire  [96:0] rsp_xbar_demux_002_src4_data;                                                                             // rsp_xbar_demux_002:src4_data -> rsp_xbar_mux_004:sink0_data
	wire  [53:0] rsp_xbar_demux_002_src4_channel;                                                                          // rsp_xbar_demux_002:src4_channel -> rsp_xbar_mux_004:sink0_channel
	wire         rsp_xbar_demux_002_src4_ready;                                                                            // rsp_xbar_mux_004:sink0_ready -> rsp_xbar_demux_002:src4_ready
	wire         rsp_xbar_demux_002_src5_endofpacket;                                                                      // rsp_xbar_demux_002:src5_endofpacket -> rsp_xbar_mux_005:sink0_endofpacket
	wire         rsp_xbar_demux_002_src5_valid;                                                                            // rsp_xbar_demux_002:src5_valid -> rsp_xbar_mux_005:sink0_valid
	wire         rsp_xbar_demux_002_src5_startofpacket;                                                                    // rsp_xbar_demux_002:src5_startofpacket -> rsp_xbar_mux_005:sink0_startofpacket
	wire  [96:0] rsp_xbar_demux_002_src5_data;                                                                             // rsp_xbar_demux_002:src5_data -> rsp_xbar_mux_005:sink0_data
	wire  [53:0] rsp_xbar_demux_002_src5_channel;                                                                          // rsp_xbar_demux_002:src5_channel -> rsp_xbar_mux_005:sink0_channel
	wire         rsp_xbar_demux_002_src5_ready;                                                                            // rsp_xbar_mux_005:sink0_ready -> rsp_xbar_demux_002:src5_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                      // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                            // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                                    // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [96:0] rsp_xbar_demux_003_src0_data;                                                                             // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire  [53:0] rsp_xbar_demux_003_src0_channel;                                                                          // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                            // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                      // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                            // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                                    // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [96:0] rsp_xbar_demux_004_src0_data;                                                                             // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire  [53:0] rsp_xbar_demux_004_src0_channel;                                                                          // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                            // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                      // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                            // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                                    // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [96:0] rsp_xbar_demux_005_src0_data;                                                                             // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire  [53:0] rsp_xbar_demux_005_src0_channel;                                                                          // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                            // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_005_src1_endofpacket;                                                                      // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire         rsp_xbar_demux_005_src1_valid;                                                                            // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_002:sink1_valid
	wire         rsp_xbar_demux_005_src1_startofpacket;                                                                    // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire  [96:0] rsp_xbar_demux_005_src1_data;                                                                             // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_002:sink1_data
	wire  [53:0] rsp_xbar_demux_005_src1_channel;                                                                          // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_002:sink1_channel
	wire         rsp_xbar_demux_005_src1_ready;                                                                            // rsp_xbar_mux_002:sink1_ready -> rsp_xbar_demux_005:src1_ready
	wire         rsp_xbar_demux_005_src2_endofpacket;                                                                      // rsp_xbar_demux_005:src2_endofpacket -> rsp_xbar_mux_004:sink1_endofpacket
	wire         rsp_xbar_demux_005_src2_valid;                                                                            // rsp_xbar_demux_005:src2_valid -> rsp_xbar_mux_004:sink1_valid
	wire         rsp_xbar_demux_005_src2_startofpacket;                                                                    // rsp_xbar_demux_005:src2_startofpacket -> rsp_xbar_mux_004:sink1_startofpacket
	wire  [96:0] rsp_xbar_demux_005_src2_data;                                                                             // rsp_xbar_demux_005:src2_data -> rsp_xbar_mux_004:sink1_data
	wire  [53:0] rsp_xbar_demux_005_src2_channel;                                                                          // rsp_xbar_demux_005:src2_channel -> rsp_xbar_mux_004:sink1_channel
	wire         rsp_xbar_demux_005_src2_ready;                                                                            // rsp_xbar_mux_004:sink1_ready -> rsp_xbar_demux_005:src2_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                      // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                            // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                                    // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [96:0] rsp_xbar_demux_006_src0_data;                                                                             // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire  [53:0] rsp_xbar_demux_006_src0_channel;                                                                          // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                            // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_006_src1_endofpacket;                                                                      // rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	wire         rsp_xbar_demux_006_src1_valid;                                                                            // rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_002:sink2_valid
	wire         rsp_xbar_demux_006_src1_startofpacket;                                                                    // rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	wire  [96:0] rsp_xbar_demux_006_src1_data;                                                                             // rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_002:sink2_data
	wire  [53:0] rsp_xbar_demux_006_src1_channel;                                                                          // rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_002:sink2_channel
	wire         rsp_xbar_demux_006_src1_ready;                                                                            // rsp_xbar_mux_002:sink2_ready -> rsp_xbar_demux_006:src1_ready
	wire         rsp_xbar_demux_006_src2_endofpacket;                                                                      // rsp_xbar_demux_006:src2_endofpacket -> rsp_xbar_mux_004:sink2_endofpacket
	wire         rsp_xbar_demux_006_src2_valid;                                                                            // rsp_xbar_demux_006:src2_valid -> rsp_xbar_mux_004:sink2_valid
	wire         rsp_xbar_demux_006_src2_startofpacket;                                                                    // rsp_xbar_demux_006:src2_startofpacket -> rsp_xbar_mux_004:sink2_startofpacket
	wire  [96:0] rsp_xbar_demux_006_src2_data;                                                                             // rsp_xbar_demux_006:src2_data -> rsp_xbar_mux_004:sink2_data
	wire  [53:0] rsp_xbar_demux_006_src2_channel;                                                                          // rsp_xbar_demux_006:src2_channel -> rsp_xbar_mux_004:sink2_channel
	wire         rsp_xbar_demux_006_src2_ready;                                                                            // rsp_xbar_mux_004:sink2_ready -> rsp_xbar_demux_006:src2_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                      // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                            // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                                    // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [96:0] rsp_xbar_demux_007_src0_data;                                                                             // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire  [53:0] rsp_xbar_demux_007_src0_channel;                                                                          // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                            // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_007_src1_endofpacket;                                                                      // rsp_xbar_demux_007:src1_endofpacket -> rsp_xbar_mux_002:sink3_endofpacket
	wire         rsp_xbar_demux_007_src1_valid;                                                                            // rsp_xbar_demux_007:src1_valid -> rsp_xbar_mux_002:sink3_valid
	wire         rsp_xbar_demux_007_src1_startofpacket;                                                                    // rsp_xbar_demux_007:src1_startofpacket -> rsp_xbar_mux_002:sink3_startofpacket
	wire  [96:0] rsp_xbar_demux_007_src1_data;                                                                             // rsp_xbar_demux_007:src1_data -> rsp_xbar_mux_002:sink3_data
	wire  [53:0] rsp_xbar_demux_007_src1_channel;                                                                          // rsp_xbar_demux_007:src1_channel -> rsp_xbar_mux_002:sink3_channel
	wire         rsp_xbar_demux_007_src1_ready;                                                                            // rsp_xbar_mux_002:sink3_ready -> rsp_xbar_demux_007:src1_ready
	wire         rsp_xbar_demux_007_src2_endofpacket;                                                                      // rsp_xbar_demux_007:src2_endofpacket -> rsp_xbar_mux_004:sink3_endofpacket
	wire         rsp_xbar_demux_007_src2_valid;                                                                            // rsp_xbar_demux_007:src2_valid -> rsp_xbar_mux_004:sink3_valid
	wire         rsp_xbar_demux_007_src2_startofpacket;                                                                    // rsp_xbar_demux_007:src2_startofpacket -> rsp_xbar_mux_004:sink3_startofpacket
	wire  [96:0] rsp_xbar_demux_007_src2_data;                                                                             // rsp_xbar_demux_007:src2_data -> rsp_xbar_mux_004:sink3_data
	wire  [53:0] rsp_xbar_demux_007_src2_channel;                                                                          // rsp_xbar_demux_007:src2_channel -> rsp_xbar_mux_004:sink3_channel
	wire         rsp_xbar_demux_007_src2_ready;                                                                            // rsp_xbar_mux_004:sink3_ready -> rsp_xbar_demux_007:src2_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                      // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                            // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                                    // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [96:0] rsp_xbar_demux_008_src0_data;                                                                             // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire  [53:0] rsp_xbar_demux_008_src0_channel;                                                                          // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                            // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_008_src1_endofpacket;                                                                      // rsp_xbar_demux_008:src1_endofpacket -> rsp_xbar_mux_002:sink4_endofpacket
	wire         rsp_xbar_demux_008_src1_valid;                                                                            // rsp_xbar_demux_008:src1_valid -> rsp_xbar_mux_002:sink4_valid
	wire         rsp_xbar_demux_008_src1_startofpacket;                                                                    // rsp_xbar_demux_008:src1_startofpacket -> rsp_xbar_mux_002:sink4_startofpacket
	wire  [96:0] rsp_xbar_demux_008_src1_data;                                                                             // rsp_xbar_demux_008:src1_data -> rsp_xbar_mux_002:sink4_data
	wire  [53:0] rsp_xbar_demux_008_src1_channel;                                                                          // rsp_xbar_demux_008:src1_channel -> rsp_xbar_mux_002:sink4_channel
	wire         rsp_xbar_demux_008_src1_ready;                                                                            // rsp_xbar_mux_002:sink4_ready -> rsp_xbar_demux_008:src1_ready
	wire         rsp_xbar_demux_008_src2_endofpacket;                                                                      // rsp_xbar_demux_008:src2_endofpacket -> rsp_xbar_mux_004:sink4_endofpacket
	wire         rsp_xbar_demux_008_src2_valid;                                                                            // rsp_xbar_demux_008:src2_valid -> rsp_xbar_mux_004:sink4_valid
	wire         rsp_xbar_demux_008_src2_startofpacket;                                                                    // rsp_xbar_demux_008:src2_startofpacket -> rsp_xbar_mux_004:sink4_startofpacket
	wire  [96:0] rsp_xbar_demux_008_src2_data;                                                                             // rsp_xbar_demux_008:src2_data -> rsp_xbar_mux_004:sink4_data
	wire  [53:0] rsp_xbar_demux_008_src2_channel;                                                                          // rsp_xbar_demux_008:src2_channel -> rsp_xbar_mux_004:sink4_channel
	wire         rsp_xbar_demux_008_src2_ready;                                                                            // rsp_xbar_mux_004:sink4_ready -> rsp_xbar_demux_008:src2_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                                      // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                            // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                                    // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [96:0] rsp_xbar_demux_009_src0_data;                                                                             // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire  [53:0] rsp_xbar_demux_009_src0_channel;                                                                          // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                            // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_009_src1_endofpacket;                                                                      // rsp_xbar_demux_009:src1_endofpacket -> rsp_xbar_mux_002:sink5_endofpacket
	wire         rsp_xbar_demux_009_src1_valid;                                                                            // rsp_xbar_demux_009:src1_valid -> rsp_xbar_mux_002:sink5_valid
	wire         rsp_xbar_demux_009_src1_startofpacket;                                                                    // rsp_xbar_demux_009:src1_startofpacket -> rsp_xbar_mux_002:sink5_startofpacket
	wire  [96:0] rsp_xbar_demux_009_src1_data;                                                                             // rsp_xbar_demux_009:src1_data -> rsp_xbar_mux_002:sink5_data
	wire  [53:0] rsp_xbar_demux_009_src1_channel;                                                                          // rsp_xbar_demux_009:src1_channel -> rsp_xbar_mux_002:sink5_channel
	wire         rsp_xbar_demux_009_src1_ready;                                                                            // rsp_xbar_mux_002:sink5_ready -> rsp_xbar_demux_009:src1_ready
	wire         rsp_xbar_demux_009_src2_endofpacket;                                                                      // rsp_xbar_demux_009:src2_endofpacket -> rsp_xbar_mux_004:sink5_endofpacket
	wire         rsp_xbar_demux_009_src2_valid;                                                                            // rsp_xbar_demux_009:src2_valid -> rsp_xbar_mux_004:sink5_valid
	wire         rsp_xbar_demux_009_src2_startofpacket;                                                                    // rsp_xbar_demux_009:src2_startofpacket -> rsp_xbar_mux_004:sink5_startofpacket
	wire  [96:0] rsp_xbar_demux_009_src2_data;                                                                             // rsp_xbar_demux_009:src2_data -> rsp_xbar_mux_004:sink5_data
	wire  [53:0] rsp_xbar_demux_009_src2_channel;                                                                          // rsp_xbar_demux_009:src2_channel -> rsp_xbar_mux_004:sink5_channel
	wire         rsp_xbar_demux_009_src2_ready;                                                                            // rsp_xbar_mux_004:sink5_ready -> rsp_xbar_demux_009:src2_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                                      // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                                            // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                                    // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [96:0] rsp_xbar_demux_010_src0_data;                                                                             // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire  [53:0] rsp_xbar_demux_010_src0_channel;                                                                          // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                                            // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire         rsp_xbar_demux_010_src1_endofpacket;                                                                      // rsp_xbar_demux_010:src1_endofpacket -> rsp_xbar_mux_002:sink6_endofpacket
	wire         rsp_xbar_demux_010_src1_valid;                                                                            // rsp_xbar_demux_010:src1_valid -> rsp_xbar_mux_002:sink6_valid
	wire         rsp_xbar_demux_010_src1_startofpacket;                                                                    // rsp_xbar_demux_010:src1_startofpacket -> rsp_xbar_mux_002:sink6_startofpacket
	wire  [96:0] rsp_xbar_demux_010_src1_data;                                                                             // rsp_xbar_demux_010:src1_data -> rsp_xbar_mux_002:sink6_data
	wire  [53:0] rsp_xbar_demux_010_src1_channel;                                                                          // rsp_xbar_demux_010:src1_channel -> rsp_xbar_mux_002:sink6_channel
	wire         rsp_xbar_demux_010_src1_ready;                                                                            // rsp_xbar_mux_002:sink6_ready -> rsp_xbar_demux_010:src1_ready
	wire         rsp_xbar_demux_010_src2_endofpacket;                                                                      // rsp_xbar_demux_010:src2_endofpacket -> rsp_xbar_mux_004:sink6_endofpacket
	wire         rsp_xbar_demux_010_src2_valid;                                                                            // rsp_xbar_demux_010:src2_valid -> rsp_xbar_mux_004:sink6_valid
	wire         rsp_xbar_demux_010_src2_startofpacket;                                                                    // rsp_xbar_demux_010:src2_startofpacket -> rsp_xbar_mux_004:sink6_startofpacket
	wire  [96:0] rsp_xbar_demux_010_src2_data;                                                                             // rsp_xbar_demux_010:src2_data -> rsp_xbar_mux_004:sink6_data
	wire  [53:0] rsp_xbar_demux_010_src2_channel;                                                                          // rsp_xbar_demux_010:src2_channel -> rsp_xbar_mux_004:sink6_channel
	wire         rsp_xbar_demux_010_src2_ready;                                                                            // rsp_xbar_mux_004:sink6_ready -> rsp_xbar_demux_010:src2_ready
	wire         rsp_xbar_demux_011_src0_endofpacket;                                                                      // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire         rsp_xbar_demux_011_src0_valid;                                                                            // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire         rsp_xbar_demux_011_src0_startofpacket;                                                                    // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [96:0] rsp_xbar_demux_011_src0_data;                                                                             // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire  [53:0] rsp_xbar_demux_011_src0_channel;                                                                          // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire         rsp_xbar_demux_011_src0_ready;                                                                            // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire         rsp_xbar_demux_012_src0_endofpacket;                                                                      // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire         rsp_xbar_demux_012_src0_valid;                                                                            // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire         rsp_xbar_demux_012_src0_startofpacket;                                                                    // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [96:0] rsp_xbar_demux_012_src0_data;                                                                             // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire  [53:0] rsp_xbar_demux_012_src0_channel;                                                                          // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire         rsp_xbar_demux_012_src0_ready;                                                                            // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire         rsp_xbar_demux_013_src0_endofpacket;                                                                      // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire         rsp_xbar_demux_013_src0_valid;                                                                            // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire         rsp_xbar_demux_013_src0_startofpacket;                                                                    // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [96:0] rsp_xbar_demux_013_src0_data;                                                                             // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire  [53:0] rsp_xbar_demux_013_src0_channel;                                                                          // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire         rsp_xbar_demux_013_src0_ready;                                                                            // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire         rsp_xbar_demux_014_src0_endofpacket;                                                                      // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire         rsp_xbar_demux_014_src0_valid;                                                                            // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	wire         rsp_xbar_demux_014_src0_startofpacket;                                                                    // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [96:0] rsp_xbar_demux_014_src0_data;                                                                             // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	wire  [53:0] rsp_xbar_demux_014_src0_channel;                                                                          // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	wire         rsp_xbar_demux_014_src0_ready;                                                                            // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire         rsp_xbar_demux_015_src0_endofpacket;                                                                      // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire         rsp_xbar_demux_015_src0_valid;                                                                            // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire         rsp_xbar_demux_015_src0_startofpacket;                                                                    // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [96:0] rsp_xbar_demux_015_src0_data;                                                                             // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire  [53:0] rsp_xbar_demux_015_src0_channel;                                                                          // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire         rsp_xbar_demux_015_src0_ready;                                                                            // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire         rsp_xbar_demux_016_src0_endofpacket;                                                                      // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire         rsp_xbar_demux_016_src0_valid;                                                                            // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	wire         rsp_xbar_demux_016_src0_startofpacket;                                                                    // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [96:0] rsp_xbar_demux_016_src0_data;                                                                             // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	wire  [53:0] rsp_xbar_demux_016_src0_channel;                                                                          // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	wire         rsp_xbar_demux_016_src0_ready;                                                                            // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire         rsp_xbar_demux_017_src0_endofpacket;                                                                      // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire         rsp_xbar_demux_017_src0_valid;                                                                            // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_001:sink17_valid
	wire         rsp_xbar_demux_017_src0_startofpacket;                                                                    // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [96:0] rsp_xbar_demux_017_src0_data;                                                                             // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_001:sink17_data
	wire  [53:0] rsp_xbar_demux_017_src0_channel;                                                                          // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_001:sink17_channel
	wire         rsp_xbar_demux_017_src0_ready;                                                                            // rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire         rsp_xbar_demux_018_src0_endofpacket;                                                                      // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire         rsp_xbar_demux_018_src0_valid;                                                                            // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_001:sink18_valid
	wire         rsp_xbar_demux_018_src0_startofpacket;                                                                    // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [96:0] rsp_xbar_demux_018_src0_data;                                                                             // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_001:sink18_data
	wire  [53:0] rsp_xbar_demux_018_src0_channel;                                                                          // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_001:sink18_channel
	wire         rsp_xbar_demux_018_src0_ready;                                                                            // rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire         rsp_xbar_demux_019_src0_endofpacket;                                                                      // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	wire         rsp_xbar_demux_019_src0_valid;                                                                            // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_001:sink19_valid
	wire         rsp_xbar_demux_019_src0_startofpacket;                                                                    // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	wire  [96:0] rsp_xbar_demux_019_src0_data;                                                                             // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_001:sink19_data
	wire  [53:0] rsp_xbar_demux_019_src0_channel;                                                                          // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_001:sink19_channel
	wire         rsp_xbar_demux_019_src0_ready;                                                                            // rsp_xbar_mux_001:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire         rsp_xbar_demux_019_src1_endofpacket;                                                                      // rsp_xbar_demux_019:src1_endofpacket -> rsp_xbar_mux_002:sink7_endofpacket
	wire         rsp_xbar_demux_019_src1_valid;                                                                            // rsp_xbar_demux_019:src1_valid -> rsp_xbar_mux_002:sink7_valid
	wire         rsp_xbar_demux_019_src1_startofpacket;                                                                    // rsp_xbar_demux_019:src1_startofpacket -> rsp_xbar_mux_002:sink7_startofpacket
	wire  [96:0] rsp_xbar_demux_019_src1_data;                                                                             // rsp_xbar_demux_019:src1_data -> rsp_xbar_mux_002:sink7_data
	wire  [53:0] rsp_xbar_demux_019_src1_channel;                                                                          // rsp_xbar_demux_019:src1_channel -> rsp_xbar_mux_002:sink7_channel
	wire         rsp_xbar_demux_019_src1_ready;                                                                            // rsp_xbar_mux_002:sink7_ready -> rsp_xbar_demux_019:src1_ready
	wire         rsp_xbar_demux_019_src2_endofpacket;                                                                      // rsp_xbar_demux_019:src2_endofpacket -> rsp_xbar_mux_004:sink7_endofpacket
	wire         rsp_xbar_demux_019_src2_valid;                                                                            // rsp_xbar_demux_019:src2_valid -> rsp_xbar_mux_004:sink7_valid
	wire         rsp_xbar_demux_019_src2_startofpacket;                                                                    // rsp_xbar_demux_019:src2_startofpacket -> rsp_xbar_mux_004:sink7_startofpacket
	wire  [96:0] rsp_xbar_demux_019_src2_data;                                                                             // rsp_xbar_demux_019:src2_data -> rsp_xbar_mux_004:sink7_data
	wire  [53:0] rsp_xbar_demux_019_src2_channel;                                                                          // rsp_xbar_demux_019:src2_channel -> rsp_xbar_mux_004:sink7_channel
	wire         rsp_xbar_demux_019_src2_ready;                                                                            // rsp_xbar_mux_004:sink7_ready -> rsp_xbar_demux_019:src2_ready
	wire         rsp_xbar_demux_020_src0_endofpacket;                                                                      // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_001:sink20_endofpacket
	wire         rsp_xbar_demux_020_src0_valid;                                                                            // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_001:sink20_valid
	wire         rsp_xbar_demux_020_src0_startofpacket;                                                                    // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_001:sink20_startofpacket
	wire  [96:0] rsp_xbar_demux_020_src0_data;                                                                             // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_001:sink20_data
	wire  [53:0] rsp_xbar_demux_020_src0_channel;                                                                          // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_001:sink20_channel
	wire         rsp_xbar_demux_020_src0_ready;                                                                            // rsp_xbar_mux_001:sink20_ready -> rsp_xbar_demux_020:src0_ready
	wire         rsp_xbar_demux_020_src1_endofpacket;                                                                      // rsp_xbar_demux_020:src1_endofpacket -> rsp_xbar_mux_002:sink8_endofpacket
	wire         rsp_xbar_demux_020_src1_valid;                                                                            // rsp_xbar_demux_020:src1_valid -> rsp_xbar_mux_002:sink8_valid
	wire         rsp_xbar_demux_020_src1_startofpacket;                                                                    // rsp_xbar_demux_020:src1_startofpacket -> rsp_xbar_mux_002:sink8_startofpacket
	wire  [96:0] rsp_xbar_demux_020_src1_data;                                                                             // rsp_xbar_demux_020:src1_data -> rsp_xbar_mux_002:sink8_data
	wire  [53:0] rsp_xbar_demux_020_src1_channel;                                                                          // rsp_xbar_demux_020:src1_channel -> rsp_xbar_mux_002:sink8_channel
	wire         rsp_xbar_demux_020_src1_ready;                                                                            // rsp_xbar_mux_002:sink8_ready -> rsp_xbar_demux_020:src1_ready
	wire         rsp_xbar_demux_020_src2_endofpacket;                                                                      // rsp_xbar_demux_020:src2_endofpacket -> rsp_xbar_mux_004:sink8_endofpacket
	wire         rsp_xbar_demux_020_src2_valid;                                                                            // rsp_xbar_demux_020:src2_valid -> rsp_xbar_mux_004:sink8_valid
	wire         rsp_xbar_demux_020_src2_startofpacket;                                                                    // rsp_xbar_demux_020:src2_startofpacket -> rsp_xbar_mux_004:sink8_startofpacket
	wire  [96:0] rsp_xbar_demux_020_src2_data;                                                                             // rsp_xbar_demux_020:src2_data -> rsp_xbar_mux_004:sink8_data
	wire  [53:0] rsp_xbar_demux_020_src2_channel;                                                                          // rsp_xbar_demux_020:src2_channel -> rsp_xbar_mux_004:sink8_channel
	wire         rsp_xbar_demux_020_src2_ready;                                                                            // rsp_xbar_mux_004:sink8_ready -> rsp_xbar_demux_020:src2_ready
	wire         rsp_xbar_demux_021_src0_endofpacket;                                                                      // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_001:sink21_endofpacket
	wire         rsp_xbar_demux_021_src0_valid;                                                                            // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_001:sink21_valid
	wire         rsp_xbar_demux_021_src0_startofpacket;                                                                    // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_001:sink21_startofpacket
	wire  [96:0] rsp_xbar_demux_021_src0_data;                                                                             // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_001:sink21_data
	wire  [53:0] rsp_xbar_demux_021_src0_channel;                                                                          // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_001:sink21_channel
	wire         rsp_xbar_demux_021_src0_ready;                                                                            // rsp_xbar_mux_001:sink21_ready -> rsp_xbar_demux_021:src0_ready
	wire         rsp_xbar_demux_021_src1_endofpacket;                                                                      // rsp_xbar_demux_021:src1_endofpacket -> rsp_xbar_mux_002:sink9_endofpacket
	wire         rsp_xbar_demux_021_src1_valid;                                                                            // rsp_xbar_demux_021:src1_valid -> rsp_xbar_mux_002:sink9_valid
	wire         rsp_xbar_demux_021_src1_startofpacket;                                                                    // rsp_xbar_demux_021:src1_startofpacket -> rsp_xbar_mux_002:sink9_startofpacket
	wire  [96:0] rsp_xbar_demux_021_src1_data;                                                                             // rsp_xbar_demux_021:src1_data -> rsp_xbar_mux_002:sink9_data
	wire  [53:0] rsp_xbar_demux_021_src1_channel;                                                                          // rsp_xbar_demux_021:src1_channel -> rsp_xbar_mux_002:sink9_channel
	wire         rsp_xbar_demux_021_src1_ready;                                                                            // rsp_xbar_mux_002:sink9_ready -> rsp_xbar_demux_021:src1_ready
	wire         rsp_xbar_demux_021_src2_endofpacket;                                                                      // rsp_xbar_demux_021:src2_endofpacket -> rsp_xbar_mux_004:sink9_endofpacket
	wire         rsp_xbar_demux_021_src2_valid;                                                                            // rsp_xbar_demux_021:src2_valid -> rsp_xbar_mux_004:sink9_valid
	wire         rsp_xbar_demux_021_src2_startofpacket;                                                                    // rsp_xbar_demux_021:src2_startofpacket -> rsp_xbar_mux_004:sink9_startofpacket
	wire  [96:0] rsp_xbar_demux_021_src2_data;                                                                             // rsp_xbar_demux_021:src2_data -> rsp_xbar_mux_004:sink9_data
	wire  [53:0] rsp_xbar_demux_021_src2_channel;                                                                          // rsp_xbar_demux_021:src2_channel -> rsp_xbar_mux_004:sink9_channel
	wire         rsp_xbar_demux_021_src2_ready;                                                                            // rsp_xbar_mux_004:sink9_ready -> rsp_xbar_demux_021:src2_ready
	wire         rsp_xbar_demux_022_src0_endofpacket;                                                                      // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_001:sink22_endofpacket
	wire         rsp_xbar_demux_022_src0_valid;                                                                            // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_001:sink22_valid
	wire         rsp_xbar_demux_022_src0_startofpacket;                                                                    // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_001:sink22_startofpacket
	wire  [96:0] rsp_xbar_demux_022_src0_data;                                                                             // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_001:sink22_data
	wire  [53:0] rsp_xbar_demux_022_src0_channel;                                                                          // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_001:sink22_channel
	wire         rsp_xbar_demux_022_src0_ready;                                                                            // rsp_xbar_mux_001:sink22_ready -> rsp_xbar_demux_022:src0_ready
	wire         rsp_xbar_demux_022_src1_endofpacket;                                                                      // rsp_xbar_demux_022:src1_endofpacket -> rsp_xbar_mux_002:sink10_endofpacket
	wire         rsp_xbar_demux_022_src1_valid;                                                                            // rsp_xbar_demux_022:src1_valid -> rsp_xbar_mux_002:sink10_valid
	wire         rsp_xbar_demux_022_src1_startofpacket;                                                                    // rsp_xbar_demux_022:src1_startofpacket -> rsp_xbar_mux_002:sink10_startofpacket
	wire  [96:0] rsp_xbar_demux_022_src1_data;                                                                             // rsp_xbar_demux_022:src1_data -> rsp_xbar_mux_002:sink10_data
	wire  [53:0] rsp_xbar_demux_022_src1_channel;                                                                          // rsp_xbar_demux_022:src1_channel -> rsp_xbar_mux_002:sink10_channel
	wire         rsp_xbar_demux_022_src1_ready;                                                                            // rsp_xbar_mux_002:sink10_ready -> rsp_xbar_demux_022:src1_ready
	wire         rsp_xbar_demux_022_src2_endofpacket;                                                                      // rsp_xbar_demux_022:src2_endofpacket -> rsp_xbar_mux_004:sink10_endofpacket
	wire         rsp_xbar_demux_022_src2_valid;                                                                            // rsp_xbar_demux_022:src2_valid -> rsp_xbar_mux_004:sink10_valid
	wire         rsp_xbar_demux_022_src2_startofpacket;                                                                    // rsp_xbar_demux_022:src2_startofpacket -> rsp_xbar_mux_004:sink10_startofpacket
	wire  [96:0] rsp_xbar_demux_022_src2_data;                                                                             // rsp_xbar_demux_022:src2_data -> rsp_xbar_mux_004:sink10_data
	wire  [53:0] rsp_xbar_demux_022_src2_channel;                                                                          // rsp_xbar_demux_022:src2_channel -> rsp_xbar_mux_004:sink10_channel
	wire         rsp_xbar_demux_022_src2_ready;                                                                            // rsp_xbar_mux_004:sink10_ready -> rsp_xbar_demux_022:src2_ready
	wire         rsp_xbar_demux_023_src0_endofpacket;                                                                      // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_001:sink23_endofpacket
	wire         rsp_xbar_demux_023_src0_valid;                                                                            // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_001:sink23_valid
	wire         rsp_xbar_demux_023_src0_startofpacket;                                                                    // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_001:sink23_startofpacket
	wire  [96:0] rsp_xbar_demux_023_src0_data;                                                                             // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_001:sink23_data
	wire  [53:0] rsp_xbar_demux_023_src0_channel;                                                                          // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_001:sink23_channel
	wire         rsp_xbar_demux_023_src0_ready;                                                                            // rsp_xbar_mux_001:sink23_ready -> rsp_xbar_demux_023:src0_ready
	wire         rsp_xbar_demux_024_src0_endofpacket;                                                                      // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_001:sink24_endofpacket
	wire         rsp_xbar_demux_024_src0_valid;                                                                            // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_001:sink24_valid
	wire         rsp_xbar_demux_024_src0_startofpacket;                                                                    // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_001:sink24_startofpacket
	wire  [96:0] rsp_xbar_demux_024_src0_data;                                                                             // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_001:sink24_data
	wire  [53:0] rsp_xbar_demux_024_src0_channel;                                                                          // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_001:sink24_channel
	wire         rsp_xbar_demux_024_src0_ready;                                                                            // rsp_xbar_mux_001:sink24_ready -> rsp_xbar_demux_024:src0_ready
	wire         rsp_xbar_demux_025_src0_endofpacket;                                                                      // rsp_xbar_demux_025:src0_endofpacket -> rsp_xbar_mux_001:sink25_endofpacket
	wire         rsp_xbar_demux_025_src0_valid;                                                                            // rsp_xbar_demux_025:src0_valid -> rsp_xbar_mux_001:sink25_valid
	wire         rsp_xbar_demux_025_src0_startofpacket;                                                                    // rsp_xbar_demux_025:src0_startofpacket -> rsp_xbar_mux_001:sink25_startofpacket
	wire  [96:0] rsp_xbar_demux_025_src0_data;                                                                             // rsp_xbar_demux_025:src0_data -> rsp_xbar_mux_001:sink25_data
	wire  [53:0] rsp_xbar_demux_025_src0_channel;                                                                          // rsp_xbar_demux_025:src0_channel -> rsp_xbar_mux_001:sink25_channel
	wire         rsp_xbar_demux_025_src0_ready;                                                                            // rsp_xbar_mux_001:sink25_ready -> rsp_xbar_demux_025:src0_ready
	wire         rsp_xbar_demux_025_src1_endofpacket;                                                                      // rsp_xbar_demux_025:src1_endofpacket -> rsp_xbar_mux_002:sink11_endofpacket
	wire         rsp_xbar_demux_025_src1_valid;                                                                            // rsp_xbar_demux_025:src1_valid -> rsp_xbar_mux_002:sink11_valid
	wire         rsp_xbar_demux_025_src1_startofpacket;                                                                    // rsp_xbar_demux_025:src1_startofpacket -> rsp_xbar_mux_002:sink11_startofpacket
	wire  [96:0] rsp_xbar_demux_025_src1_data;                                                                             // rsp_xbar_demux_025:src1_data -> rsp_xbar_mux_002:sink11_data
	wire  [53:0] rsp_xbar_demux_025_src1_channel;                                                                          // rsp_xbar_demux_025:src1_channel -> rsp_xbar_mux_002:sink11_channel
	wire         rsp_xbar_demux_025_src1_ready;                                                                            // rsp_xbar_mux_002:sink11_ready -> rsp_xbar_demux_025:src1_ready
	wire         rsp_xbar_demux_025_src2_endofpacket;                                                                      // rsp_xbar_demux_025:src2_endofpacket -> rsp_xbar_mux_004:sink11_endofpacket
	wire         rsp_xbar_demux_025_src2_valid;                                                                            // rsp_xbar_demux_025:src2_valid -> rsp_xbar_mux_004:sink11_valid
	wire         rsp_xbar_demux_025_src2_startofpacket;                                                                    // rsp_xbar_demux_025:src2_startofpacket -> rsp_xbar_mux_004:sink11_startofpacket
	wire  [96:0] rsp_xbar_demux_025_src2_data;                                                                             // rsp_xbar_demux_025:src2_data -> rsp_xbar_mux_004:sink11_data
	wire  [53:0] rsp_xbar_demux_025_src2_channel;                                                                          // rsp_xbar_demux_025:src2_channel -> rsp_xbar_mux_004:sink11_channel
	wire         rsp_xbar_demux_025_src2_ready;                                                                            // rsp_xbar_mux_004:sink11_ready -> rsp_xbar_demux_025:src2_ready
	wire         rsp_xbar_demux_026_src0_endofpacket;                                                                      // rsp_xbar_demux_026:src0_endofpacket -> rsp_xbar_mux_002:sink12_endofpacket
	wire         rsp_xbar_demux_026_src0_valid;                                                                            // rsp_xbar_demux_026:src0_valid -> rsp_xbar_mux_002:sink12_valid
	wire         rsp_xbar_demux_026_src0_startofpacket;                                                                    // rsp_xbar_demux_026:src0_startofpacket -> rsp_xbar_mux_002:sink12_startofpacket
	wire  [96:0] rsp_xbar_demux_026_src0_data;                                                                             // rsp_xbar_demux_026:src0_data -> rsp_xbar_mux_002:sink12_data
	wire  [53:0] rsp_xbar_demux_026_src0_channel;                                                                          // rsp_xbar_demux_026:src0_channel -> rsp_xbar_mux_002:sink12_channel
	wire         rsp_xbar_demux_026_src0_ready;                                                                            // rsp_xbar_mux_002:sink12_ready -> rsp_xbar_demux_026:src0_ready
	wire         rsp_xbar_demux_026_src1_endofpacket;                                                                      // rsp_xbar_demux_026:src1_endofpacket -> rsp_xbar_mux_003:sink1_endofpacket
	wire         rsp_xbar_demux_026_src1_valid;                                                                            // rsp_xbar_demux_026:src1_valid -> rsp_xbar_mux_003:sink1_valid
	wire         rsp_xbar_demux_026_src1_startofpacket;                                                                    // rsp_xbar_demux_026:src1_startofpacket -> rsp_xbar_mux_003:sink1_startofpacket
	wire  [96:0] rsp_xbar_demux_026_src1_data;                                                                             // rsp_xbar_demux_026:src1_data -> rsp_xbar_mux_003:sink1_data
	wire  [53:0] rsp_xbar_demux_026_src1_channel;                                                                          // rsp_xbar_demux_026:src1_channel -> rsp_xbar_mux_003:sink1_channel
	wire         rsp_xbar_demux_026_src1_ready;                                                                            // rsp_xbar_mux_003:sink1_ready -> rsp_xbar_demux_026:src1_ready
	wire         rsp_xbar_demux_027_src0_endofpacket;                                                                      // rsp_xbar_demux_027:src0_endofpacket -> rsp_xbar_mux_002:sink13_endofpacket
	wire         rsp_xbar_demux_027_src0_valid;                                                                            // rsp_xbar_demux_027:src0_valid -> rsp_xbar_mux_002:sink13_valid
	wire         rsp_xbar_demux_027_src0_startofpacket;                                                                    // rsp_xbar_demux_027:src0_startofpacket -> rsp_xbar_mux_002:sink13_startofpacket
	wire  [96:0] rsp_xbar_demux_027_src0_data;                                                                             // rsp_xbar_demux_027:src0_data -> rsp_xbar_mux_002:sink13_data
	wire  [53:0] rsp_xbar_demux_027_src0_channel;                                                                          // rsp_xbar_demux_027:src0_channel -> rsp_xbar_mux_002:sink13_channel
	wire         rsp_xbar_demux_027_src0_ready;                                                                            // rsp_xbar_mux_002:sink13_ready -> rsp_xbar_demux_027:src0_ready
	wire         rsp_xbar_demux_027_src1_endofpacket;                                                                      // rsp_xbar_demux_027:src1_endofpacket -> rsp_xbar_mux_003:sink2_endofpacket
	wire         rsp_xbar_demux_027_src1_valid;                                                                            // rsp_xbar_demux_027:src1_valid -> rsp_xbar_mux_003:sink2_valid
	wire         rsp_xbar_demux_027_src1_startofpacket;                                                                    // rsp_xbar_demux_027:src1_startofpacket -> rsp_xbar_mux_003:sink2_startofpacket
	wire  [96:0] rsp_xbar_demux_027_src1_data;                                                                             // rsp_xbar_demux_027:src1_data -> rsp_xbar_mux_003:sink2_data
	wire  [53:0] rsp_xbar_demux_027_src1_channel;                                                                          // rsp_xbar_demux_027:src1_channel -> rsp_xbar_mux_003:sink2_channel
	wire         rsp_xbar_demux_027_src1_ready;                                                                            // rsp_xbar_mux_003:sink2_ready -> rsp_xbar_demux_027:src1_ready
	wire         rsp_xbar_demux_028_src0_endofpacket;                                                                      // rsp_xbar_demux_028:src0_endofpacket -> rsp_xbar_mux_002:sink14_endofpacket
	wire         rsp_xbar_demux_028_src0_valid;                                                                            // rsp_xbar_demux_028:src0_valid -> rsp_xbar_mux_002:sink14_valid
	wire         rsp_xbar_demux_028_src0_startofpacket;                                                                    // rsp_xbar_demux_028:src0_startofpacket -> rsp_xbar_mux_002:sink14_startofpacket
	wire  [96:0] rsp_xbar_demux_028_src0_data;                                                                             // rsp_xbar_demux_028:src0_data -> rsp_xbar_mux_002:sink14_data
	wire  [53:0] rsp_xbar_demux_028_src0_channel;                                                                          // rsp_xbar_demux_028:src0_channel -> rsp_xbar_mux_002:sink14_channel
	wire         rsp_xbar_demux_028_src0_ready;                                                                            // rsp_xbar_mux_002:sink14_ready -> rsp_xbar_demux_028:src0_ready
	wire         rsp_xbar_demux_029_src0_endofpacket;                                                                      // rsp_xbar_demux_029:src0_endofpacket -> rsp_xbar_mux_002:sink15_endofpacket
	wire         rsp_xbar_demux_029_src0_valid;                                                                            // rsp_xbar_demux_029:src0_valid -> rsp_xbar_mux_002:sink15_valid
	wire         rsp_xbar_demux_029_src0_startofpacket;                                                                    // rsp_xbar_demux_029:src0_startofpacket -> rsp_xbar_mux_002:sink15_startofpacket
	wire  [96:0] rsp_xbar_demux_029_src0_data;                                                                             // rsp_xbar_demux_029:src0_data -> rsp_xbar_mux_002:sink15_data
	wire  [53:0] rsp_xbar_demux_029_src0_channel;                                                                          // rsp_xbar_demux_029:src0_channel -> rsp_xbar_mux_002:sink15_channel
	wire         rsp_xbar_demux_029_src0_ready;                                                                            // rsp_xbar_mux_002:sink15_ready -> rsp_xbar_demux_029:src0_ready
	wire         rsp_xbar_demux_030_src0_endofpacket;                                                                      // rsp_xbar_demux_030:src0_endofpacket -> rsp_xbar_mux_002:sink16_endofpacket
	wire         rsp_xbar_demux_030_src0_valid;                                                                            // rsp_xbar_demux_030:src0_valid -> rsp_xbar_mux_002:sink16_valid
	wire         rsp_xbar_demux_030_src0_startofpacket;                                                                    // rsp_xbar_demux_030:src0_startofpacket -> rsp_xbar_mux_002:sink16_startofpacket
	wire  [96:0] rsp_xbar_demux_030_src0_data;                                                                             // rsp_xbar_demux_030:src0_data -> rsp_xbar_mux_002:sink16_data
	wire  [53:0] rsp_xbar_demux_030_src0_channel;                                                                          // rsp_xbar_demux_030:src0_channel -> rsp_xbar_mux_002:sink16_channel
	wire         rsp_xbar_demux_030_src0_ready;                                                                            // rsp_xbar_mux_002:sink16_ready -> rsp_xbar_demux_030:src0_ready
	wire         rsp_xbar_demux_031_src0_endofpacket;                                                                      // rsp_xbar_demux_031:src0_endofpacket -> rsp_xbar_mux_002:sink17_endofpacket
	wire         rsp_xbar_demux_031_src0_valid;                                                                            // rsp_xbar_demux_031:src0_valid -> rsp_xbar_mux_002:sink17_valid
	wire         rsp_xbar_demux_031_src0_startofpacket;                                                                    // rsp_xbar_demux_031:src0_startofpacket -> rsp_xbar_mux_002:sink17_startofpacket
	wire  [96:0] rsp_xbar_demux_031_src0_data;                                                                             // rsp_xbar_demux_031:src0_data -> rsp_xbar_mux_002:sink17_data
	wire  [53:0] rsp_xbar_demux_031_src0_channel;                                                                          // rsp_xbar_demux_031:src0_channel -> rsp_xbar_mux_002:sink17_channel
	wire         rsp_xbar_demux_031_src0_ready;                                                                            // rsp_xbar_mux_002:sink17_ready -> rsp_xbar_demux_031:src0_ready
	wire         rsp_xbar_demux_032_src0_endofpacket;                                                                      // rsp_xbar_demux_032:src0_endofpacket -> rsp_xbar_mux_002:sink18_endofpacket
	wire         rsp_xbar_demux_032_src0_valid;                                                                            // rsp_xbar_demux_032:src0_valid -> rsp_xbar_mux_002:sink18_valid
	wire         rsp_xbar_demux_032_src0_startofpacket;                                                                    // rsp_xbar_demux_032:src0_startofpacket -> rsp_xbar_mux_002:sink18_startofpacket
	wire  [96:0] rsp_xbar_demux_032_src0_data;                                                                             // rsp_xbar_demux_032:src0_data -> rsp_xbar_mux_002:sink18_data
	wire  [53:0] rsp_xbar_demux_032_src0_channel;                                                                          // rsp_xbar_demux_032:src0_channel -> rsp_xbar_mux_002:sink18_channel
	wire         rsp_xbar_demux_032_src0_ready;                                                                            // rsp_xbar_mux_002:sink18_ready -> rsp_xbar_demux_032:src0_ready
	wire         rsp_xbar_demux_033_src0_endofpacket;                                                                      // rsp_xbar_demux_033:src0_endofpacket -> rsp_xbar_mux_002:sink19_endofpacket
	wire         rsp_xbar_demux_033_src0_valid;                                                                            // rsp_xbar_demux_033:src0_valid -> rsp_xbar_mux_002:sink19_valid
	wire         rsp_xbar_demux_033_src0_startofpacket;                                                                    // rsp_xbar_demux_033:src0_startofpacket -> rsp_xbar_mux_002:sink19_startofpacket
	wire  [96:0] rsp_xbar_demux_033_src0_data;                                                                             // rsp_xbar_demux_033:src0_data -> rsp_xbar_mux_002:sink19_data
	wire  [53:0] rsp_xbar_demux_033_src0_channel;                                                                          // rsp_xbar_demux_033:src0_channel -> rsp_xbar_mux_002:sink19_channel
	wire         rsp_xbar_demux_033_src0_ready;                                                                            // rsp_xbar_mux_002:sink19_ready -> rsp_xbar_demux_033:src0_ready
	wire         rsp_xbar_demux_034_src0_endofpacket;                                                                      // rsp_xbar_demux_034:src0_endofpacket -> rsp_xbar_mux_002:sink20_endofpacket
	wire         rsp_xbar_demux_034_src0_valid;                                                                            // rsp_xbar_demux_034:src0_valid -> rsp_xbar_mux_002:sink20_valid
	wire         rsp_xbar_demux_034_src0_startofpacket;                                                                    // rsp_xbar_demux_034:src0_startofpacket -> rsp_xbar_mux_002:sink20_startofpacket
	wire  [96:0] rsp_xbar_demux_034_src0_data;                                                                             // rsp_xbar_demux_034:src0_data -> rsp_xbar_mux_002:sink20_data
	wire  [53:0] rsp_xbar_demux_034_src0_channel;                                                                          // rsp_xbar_demux_034:src0_channel -> rsp_xbar_mux_002:sink20_channel
	wire         rsp_xbar_demux_034_src0_ready;                                                                            // rsp_xbar_mux_002:sink20_ready -> rsp_xbar_demux_034:src0_ready
	wire         rsp_xbar_demux_035_src0_endofpacket;                                                                      // rsp_xbar_demux_035:src0_endofpacket -> rsp_xbar_mux_002:sink21_endofpacket
	wire         rsp_xbar_demux_035_src0_valid;                                                                            // rsp_xbar_demux_035:src0_valid -> rsp_xbar_mux_002:sink21_valid
	wire         rsp_xbar_demux_035_src0_startofpacket;                                                                    // rsp_xbar_demux_035:src0_startofpacket -> rsp_xbar_mux_002:sink21_startofpacket
	wire  [96:0] rsp_xbar_demux_035_src0_data;                                                                             // rsp_xbar_demux_035:src0_data -> rsp_xbar_mux_002:sink21_data
	wire  [53:0] rsp_xbar_demux_035_src0_channel;                                                                          // rsp_xbar_demux_035:src0_channel -> rsp_xbar_mux_002:sink21_channel
	wire         rsp_xbar_demux_035_src0_ready;                                                                            // rsp_xbar_mux_002:sink21_ready -> rsp_xbar_demux_035:src0_ready
	wire         rsp_xbar_demux_036_src0_endofpacket;                                                                      // rsp_xbar_demux_036:src0_endofpacket -> rsp_xbar_mux_002:sink22_endofpacket
	wire         rsp_xbar_demux_036_src0_valid;                                                                            // rsp_xbar_demux_036:src0_valid -> rsp_xbar_mux_002:sink22_valid
	wire         rsp_xbar_demux_036_src0_startofpacket;                                                                    // rsp_xbar_demux_036:src0_startofpacket -> rsp_xbar_mux_002:sink22_startofpacket
	wire  [96:0] rsp_xbar_demux_036_src0_data;                                                                             // rsp_xbar_demux_036:src0_data -> rsp_xbar_mux_002:sink22_data
	wire  [53:0] rsp_xbar_demux_036_src0_channel;                                                                          // rsp_xbar_demux_036:src0_channel -> rsp_xbar_mux_002:sink22_channel
	wire         rsp_xbar_demux_036_src0_ready;                                                                            // rsp_xbar_mux_002:sink22_ready -> rsp_xbar_demux_036:src0_ready
	wire         rsp_xbar_demux_037_src0_endofpacket;                                                                      // rsp_xbar_demux_037:src0_endofpacket -> rsp_xbar_mux_002:sink23_endofpacket
	wire         rsp_xbar_demux_037_src0_valid;                                                                            // rsp_xbar_demux_037:src0_valid -> rsp_xbar_mux_002:sink23_valid
	wire         rsp_xbar_demux_037_src0_startofpacket;                                                                    // rsp_xbar_demux_037:src0_startofpacket -> rsp_xbar_mux_002:sink23_startofpacket
	wire  [96:0] rsp_xbar_demux_037_src0_data;                                                                             // rsp_xbar_demux_037:src0_data -> rsp_xbar_mux_002:sink23_data
	wire  [53:0] rsp_xbar_demux_037_src0_channel;                                                                          // rsp_xbar_demux_037:src0_channel -> rsp_xbar_mux_002:sink23_channel
	wire         rsp_xbar_demux_037_src0_ready;                                                                            // rsp_xbar_mux_002:sink23_ready -> rsp_xbar_demux_037:src0_ready
	wire         rsp_xbar_demux_038_src0_endofpacket;                                                                      // rsp_xbar_demux_038:src0_endofpacket -> rsp_xbar_mux_002:sink24_endofpacket
	wire         rsp_xbar_demux_038_src0_valid;                                                                            // rsp_xbar_demux_038:src0_valid -> rsp_xbar_mux_002:sink24_valid
	wire         rsp_xbar_demux_038_src0_startofpacket;                                                                    // rsp_xbar_demux_038:src0_startofpacket -> rsp_xbar_mux_002:sink24_startofpacket
	wire  [96:0] rsp_xbar_demux_038_src0_data;                                                                             // rsp_xbar_demux_038:src0_data -> rsp_xbar_mux_002:sink24_data
	wire  [53:0] rsp_xbar_demux_038_src0_channel;                                                                          // rsp_xbar_demux_038:src0_channel -> rsp_xbar_mux_002:sink24_channel
	wire         rsp_xbar_demux_038_src0_ready;                                                                            // rsp_xbar_mux_002:sink24_ready -> rsp_xbar_demux_038:src0_ready
	wire         rsp_xbar_demux_039_src0_endofpacket;                                                                      // rsp_xbar_demux_039:src0_endofpacket -> rsp_xbar_mux_002:sink25_endofpacket
	wire         rsp_xbar_demux_039_src0_valid;                                                                            // rsp_xbar_demux_039:src0_valid -> rsp_xbar_mux_002:sink25_valid
	wire         rsp_xbar_demux_039_src0_startofpacket;                                                                    // rsp_xbar_demux_039:src0_startofpacket -> rsp_xbar_mux_002:sink25_startofpacket
	wire  [96:0] rsp_xbar_demux_039_src0_data;                                                                             // rsp_xbar_demux_039:src0_data -> rsp_xbar_mux_002:sink25_data
	wire  [53:0] rsp_xbar_demux_039_src0_channel;                                                                          // rsp_xbar_demux_039:src0_channel -> rsp_xbar_mux_002:sink25_channel
	wire         rsp_xbar_demux_039_src0_ready;                                                                            // rsp_xbar_mux_002:sink25_ready -> rsp_xbar_demux_039:src0_ready
	wire         rsp_xbar_demux_040_src0_endofpacket;                                                                      // rsp_xbar_demux_040:src0_endofpacket -> rsp_xbar_mux_004:sink12_endofpacket
	wire         rsp_xbar_demux_040_src0_valid;                                                                            // rsp_xbar_demux_040:src0_valid -> rsp_xbar_mux_004:sink12_valid
	wire         rsp_xbar_demux_040_src0_startofpacket;                                                                    // rsp_xbar_demux_040:src0_startofpacket -> rsp_xbar_mux_004:sink12_startofpacket
	wire  [96:0] rsp_xbar_demux_040_src0_data;                                                                             // rsp_xbar_demux_040:src0_data -> rsp_xbar_mux_004:sink12_data
	wire  [53:0] rsp_xbar_demux_040_src0_channel;                                                                          // rsp_xbar_demux_040:src0_channel -> rsp_xbar_mux_004:sink12_channel
	wire         rsp_xbar_demux_040_src0_ready;                                                                            // rsp_xbar_mux_004:sink12_ready -> rsp_xbar_demux_040:src0_ready
	wire         rsp_xbar_demux_040_src1_endofpacket;                                                                      // rsp_xbar_demux_040:src1_endofpacket -> rsp_xbar_mux_005:sink1_endofpacket
	wire         rsp_xbar_demux_040_src1_valid;                                                                            // rsp_xbar_demux_040:src1_valid -> rsp_xbar_mux_005:sink1_valid
	wire         rsp_xbar_demux_040_src1_startofpacket;                                                                    // rsp_xbar_demux_040:src1_startofpacket -> rsp_xbar_mux_005:sink1_startofpacket
	wire  [96:0] rsp_xbar_demux_040_src1_data;                                                                             // rsp_xbar_demux_040:src1_data -> rsp_xbar_mux_005:sink1_data
	wire  [53:0] rsp_xbar_demux_040_src1_channel;                                                                          // rsp_xbar_demux_040:src1_channel -> rsp_xbar_mux_005:sink1_channel
	wire         rsp_xbar_demux_040_src1_ready;                                                                            // rsp_xbar_mux_005:sink1_ready -> rsp_xbar_demux_040:src1_ready
	wire         rsp_xbar_demux_041_src0_endofpacket;                                                                      // rsp_xbar_demux_041:src0_endofpacket -> rsp_xbar_mux_004:sink13_endofpacket
	wire         rsp_xbar_demux_041_src0_valid;                                                                            // rsp_xbar_demux_041:src0_valid -> rsp_xbar_mux_004:sink13_valid
	wire         rsp_xbar_demux_041_src0_startofpacket;                                                                    // rsp_xbar_demux_041:src0_startofpacket -> rsp_xbar_mux_004:sink13_startofpacket
	wire  [96:0] rsp_xbar_demux_041_src0_data;                                                                             // rsp_xbar_demux_041:src0_data -> rsp_xbar_mux_004:sink13_data
	wire  [53:0] rsp_xbar_demux_041_src0_channel;                                                                          // rsp_xbar_demux_041:src0_channel -> rsp_xbar_mux_004:sink13_channel
	wire         rsp_xbar_demux_041_src0_ready;                                                                            // rsp_xbar_mux_004:sink13_ready -> rsp_xbar_demux_041:src0_ready
	wire         rsp_xbar_demux_041_src1_endofpacket;                                                                      // rsp_xbar_demux_041:src1_endofpacket -> rsp_xbar_mux_005:sink2_endofpacket
	wire         rsp_xbar_demux_041_src1_valid;                                                                            // rsp_xbar_demux_041:src1_valid -> rsp_xbar_mux_005:sink2_valid
	wire         rsp_xbar_demux_041_src1_startofpacket;                                                                    // rsp_xbar_demux_041:src1_startofpacket -> rsp_xbar_mux_005:sink2_startofpacket
	wire  [96:0] rsp_xbar_demux_041_src1_data;                                                                             // rsp_xbar_demux_041:src1_data -> rsp_xbar_mux_005:sink2_data
	wire  [53:0] rsp_xbar_demux_041_src1_channel;                                                                          // rsp_xbar_demux_041:src1_channel -> rsp_xbar_mux_005:sink2_channel
	wire         rsp_xbar_demux_041_src1_ready;                                                                            // rsp_xbar_mux_005:sink2_ready -> rsp_xbar_demux_041:src1_ready
	wire         rsp_xbar_demux_042_src0_endofpacket;                                                                      // rsp_xbar_demux_042:src0_endofpacket -> rsp_xbar_mux_004:sink14_endofpacket
	wire         rsp_xbar_demux_042_src0_valid;                                                                            // rsp_xbar_demux_042:src0_valid -> rsp_xbar_mux_004:sink14_valid
	wire         rsp_xbar_demux_042_src0_startofpacket;                                                                    // rsp_xbar_demux_042:src0_startofpacket -> rsp_xbar_mux_004:sink14_startofpacket
	wire  [96:0] rsp_xbar_demux_042_src0_data;                                                                             // rsp_xbar_demux_042:src0_data -> rsp_xbar_mux_004:sink14_data
	wire  [53:0] rsp_xbar_demux_042_src0_channel;                                                                          // rsp_xbar_demux_042:src0_channel -> rsp_xbar_mux_004:sink14_channel
	wire         rsp_xbar_demux_042_src0_ready;                                                                            // rsp_xbar_mux_004:sink14_ready -> rsp_xbar_demux_042:src0_ready
	wire         rsp_xbar_demux_043_src0_endofpacket;                                                                      // rsp_xbar_demux_043:src0_endofpacket -> rsp_xbar_mux_004:sink15_endofpacket
	wire         rsp_xbar_demux_043_src0_valid;                                                                            // rsp_xbar_demux_043:src0_valid -> rsp_xbar_mux_004:sink15_valid
	wire         rsp_xbar_demux_043_src0_startofpacket;                                                                    // rsp_xbar_demux_043:src0_startofpacket -> rsp_xbar_mux_004:sink15_startofpacket
	wire  [96:0] rsp_xbar_demux_043_src0_data;                                                                             // rsp_xbar_demux_043:src0_data -> rsp_xbar_mux_004:sink15_data
	wire  [53:0] rsp_xbar_demux_043_src0_channel;                                                                          // rsp_xbar_demux_043:src0_channel -> rsp_xbar_mux_004:sink15_channel
	wire         rsp_xbar_demux_043_src0_ready;                                                                            // rsp_xbar_mux_004:sink15_ready -> rsp_xbar_demux_043:src0_ready
	wire         rsp_xbar_demux_044_src0_endofpacket;                                                                      // rsp_xbar_demux_044:src0_endofpacket -> rsp_xbar_mux_004:sink16_endofpacket
	wire         rsp_xbar_demux_044_src0_valid;                                                                            // rsp_xbar_demux_044:src0_valid -> rsp_xbar_mux_004:sink16_valid
	wire         rsp_xbar_demux_044_src0_startofpacket;                                                                    // rsp_xbar_demux_044:src0_startofpacket -> rsp_xbar_mux_004:sink16_startofpacket
	wire  [96:0] rsp_xbar_demux_044_src0_data;                                                                             // rsp_xbar_demux_044:src0_data -> rsp_xbar_mux_004:sink16_data
	wire  [53:0] rsp_xbar_demux_044_src0_channel;                                                                          // rsp_xbar_demux_044:src0_channel -> rsp_xbar_mux_004:sink16_channel
	wire         rsp_xbar_demux_044_src0_ready;                                                                            // rsp_xbar_mux_004:sink16_ready -> rsp_xbar_demux_044:src0_ready
	wire         rsp_xbar_demux_045_src0_endofpacket;                                                                      // rsp_xbar_demux_045:src0_endofpacket -> rsp_xbar_mux_004:sink17_endofpacket
	wire         rsp_xbar_demux_045_src0_valid;                                                                            // rsp_xbar_demux_045:src0_valid -> rsp_xbar_mux_004:sink17_valid
	wire         rsp_xbar_demux_045_src0_startofpacket;                                                                    // rsp_xbar_demux_045:src0_startofpacket -> rsp_xbar_mux_004:sink17_startofpacket
	wire  [96:0] rsp_xbar_demux_045_src0_data;                                                                             // rsp_xbar_demux_045:src0_data -> rsp_xbar_mux_004:sink17_data
	wire  [53:0] rsp_xbar_demux_045_src0_channel;                                                                          // rsp_xbar_demux_045:src0_channel -> rsp_xbar_mux_004:sink17_channel
	wire         rsp_xbar_demux_045_src0_ready;                                                                            // rsp_xbar_mux_004:sink17_ready -> rsp_xbar_demux_045:src0_ready
	wire         rsp_xbar_demux_046_src0_endofpacket;                                                                      // rsp_xbar_demux_046:src0_endofpacket -> rsp_xbar_mux_004:sink18_endofpacket
	wire         rsp_xbar_demux_046_src0_valid;                                                                            // rsp_xbar_demux_046:src0_valid -> rsp_xbar_mux_004:sink18_valid
	wire         rsp_xbar_demux_046_src0_startofpacket;                                                                    // rsp_xbar_demux_046:src0_startofpacket -> rsp_xbar_mux_004:sink18_startofpacket
	wire  [96:0] rsp_xbar_demux_046_src0_data;                                                                             // rsp_xbar_demux_046:src0_data -> rsp_xbar_mux_004:sink18_data
	wire  [53:0] rsp_xbar_demux_046_src0_channel;                                                                          // rsp_xbar_demux_046:src0_channel -> rsp_xbar_mux_004:sink18_channel
	wire         rsp_xbar_demux_046_src0_ready;                                                                            // rsp_xbar_mux_004:sink18_ready -> rsp_xbar_demux_046:src0_ready
	wire         rsp_xbar_demux_047_src0_endofpacket;                                                                      // rsp_xbar_demux_047:src0_endofpacket -> rsp_xbar_mux_004:sink19_endofpacket
	wire         rsp_xbar_demux_047_src0_valid;                                                                            // rsp_xbar_demux_047:src0_valid -> rsp_xbar_mux_004:sink19_valid
	wire         rsp_xbar_demux_047_src0_startofpacket;                                                                    // rsp_xbar_demux_047:src0_startofpacket -> rsp_xbar_mux_004:sink19_startofpacket
	wire  [96:0] rsp_xbar_demux_047_src0_data;                                                                             // rsp_xbar_demux_047:src0_data -> rsp_xbar_mux_004:sink19_data
	wire  [53:0] rsp_xbar_demux_047_src0_channel;                                                                          // rsp_xbar_demux_047:src0_channel -> rsp_xbar_mux_004:sink19_channel
	wire         rsp_xbar_demux_047_src0_ready;                                                                            // rsp_xbar_mux_004:sink19_ready -> rsp_xbar_demux_047:src0_ready
	wire         rsp_xbar_demux_048_src0_endofpacket;                                                                      // rsp_xbar_demux_048:src0_endofpacket -> rsp_xbar_mux_004:sink20_endofpacket
	wire         rsp_xbar_demux_048_src0_valid;                                                                            // rsp_xbar_demux_048:src0_valid -> rsp_xbar_mux_004:sink20_valid
	wire         rsp_xbar_demux_048_src0_startofpacket;                                                                    // rsp_xbar_demux_048:src0_startofpacket -> rsp_xbar_mux_004:sink20_startofpacket
	wire  [96:0] rsp_xbar_demux_048_src0_data;                                                                             // rsp_xbar_demux_048:src0_data -> rsp_xbar_mux_004:sink20_data
	wire  [53:0] rsp_xbar_demux_048_src0_channel;                                                                          // rsp_xbar_demux_048:src0_channel -> rsp_xbar_mux_004:sink20_channel
	wire         rsp_xbar_demux_048_src0_ready;                                                                            // rsp_xbar_mux_004:sink20_ready -> rsp_xbar_demux_048:src0_ready
	wire         rsp_xbar_demux_049_src0_endofpacket;                                                                      // rsp_xbar_demux_049:src0_endofpacket -> rsp_xbar_mux_004:sink21_endofpacket
	wire         rsp_xbar_demux_049_src0_valid;                                                                            // rsp_xbar_demux_049:src0_valid -> rsp_xbar_mux_004:sink21_valid
	wire         rsp_xbar_demux_049_src0_startofpacket;                                                                    // rsp_xbar_demux_049:src0_startofpacket -> rsp_xbar_mux_004:sink21_startofpacket
	wire  [96:0] rsp_xbar_demux_049_src0_data;                                                                             // rsp_xbar_demux_049:src0_data -> rsp_xbar_mux_004:sink21_data
	wire  [53:0] rsp_xbar_demux_049_src0_channel;                                                                          // rsp_xbar_demux_049:src0_channel -> rsp_xbar_mux_004:sink21_channel
	wire         rsp_xbar_demux_049_src0_ready;                                                                            // rsp_xbar_mux_004:sink21_ready -> rsp_xbar_demux_049:src0_ready
	wire         rsp_xbar_demux_050_src0_endofpacket;                                                                      // rsp_xbar_demux_050:src0_endofpacket -> rsp_xbar_mux_004:sink22_endofpacket
	wire         rsp_xbar_demux_050_src0_valid;                                                                            // rsp_xbar_demux_050:src0_valid -> rsp_xbar_mux_004:sink22_valid
	wire         rsp_xbar_demux_050_src0_startofpacket;                                                                    // rsp_xbar_demux_050:src0_startofpacket -> rsp_xbar_mux_004:sink22_startofpacket
	wire  [96:0] rsp_xbar_demux_050_src0_data;                                                                             // rsp_xbar_demux_050:src0_data -> rsp_xbar_mux_004:sink22_data
	wire  [53:0] rsp_xbar_demux_050_src0_channel;                                                                          // rsp_xbar_demux_050:src0_channel -> rsp_xbar_mux_004:sink22_channel
	wire         rsp_xbar_demux_050_src0_ready;                                                                            // rsp_xbar_mux_004:sink22_ready -> rsp_xbar_demux_050:src0_ready
	wire         rsp_xbar_demux_051_src0_endofpacket;                                                                      // rsp_xbar_demux_051:src0_endofpacket -> rsp_xbar_mux_004:sink23_endofpacket
	wire         rsp_xbar_demux_051_src0_valid;                                                                            // rsp_xbar_demux_051:src0_valid -> rsp_xbar_mux_004:sink23_valid
	wire         rsp_xbar_demux_051_src0_startofpacket;                                                                    // rsp_xbar_demux_051:src0_startofpacket -> rsp_xbar_mux_004:sink23_startofpacket
	wire  [96:0] rsp_xbar_demux_051_src0_data;                                                                             // rsp_xbar_demux_051:src0_data -> rsp_xbar_mux_004:sink23_data
	wire  [53:0] rsp_xbar_demux_051_src0_channel;                                                                          // rsp_xbar_demux_051:src0_channel -> rsp_xbar_mux_004:sink23_channel
	wire         rsp_xbar_demux_051_src0_ready;                                                                            // rsp_xbar_mux_004:sink23_ready -> rsp_xbar_demux_051:src0_ready
	wire         rsp_xbar_demux_052_src0_endofpacket;                                                                      // rsp_xbar_demux_052:src0_endofpacket -> rsp_xbar_mux_004:sink24_endofpacket
	wire         rsp_xbar_demux_052_src0_valid;                                                                            // rsp_xbar_demux_052:src0_valid -> rsp_xbar_mux_004:sink24_valid
	wire         rsp_xbar_demux_052_src0_startofpacket;                                                                    // rsp_xbar_demux_052:src0_startofpacket -> rsp_xbar_mux_004:sink24_startofpacket
	wire  [96:0] rsp_xbar_demux_052_src0_data;                                                                             // rsp_xbar_demux_052:src0_data -> rsp_xbar_mux_004:sink24_data
	wire  [53:0] rsp_xbar_demux_052_src0_channel;                                                                          // rsp_xbar_demux_052:src0_channel -> rsp_xbar_mux_004:sink24_channel
	wire         rsp_xbar_demux_052_src0_ready;                                                                            // rsp_xbar_mux_004:sink24_ready -> rsp_xbar_demux_052:src0_ready
	wire         rsp_xbar_demux_053_src0_endofpacket;                                                                      // rsp_xbar_demux_053:src0_endofpacket -> rsp_xbar_mux_004:sink25_endofpacket
	wire         rsp_xbar_demux_053_src0_valid;                                                                            // rsp_xbar_demux_053:src0_valid -> rsp_xbar_mux_004:sink25_valid
	wire         rsp_xbar_demux_053_src0_startofpacket;                                                                    // rsp_xbar_demux_053:src0_startofpacket -> rsp_xbar_mux_004:sink25_startofpacket
	wire  [96:0] rsp_xbar_demux_053_src0_data;                                                                             // rsp_xbar_demux_053:src0_data -> rsp_xbar_mux_004:sink25_data
	wire  [53:0] rsp_xbar_demux_053_src0_channel;                                                                          // rsp_xbar_demux_053:src0_channel -> rsp_xbar_mux_004:sink25_channel
	wire         rsp_xbar_demux_053_src0_ready;                                                                            // rsp_xbar_mux_004:sink25_ready -> rsp_xbar_demux_053:src0_ready
	wire         addr_router_src_endofpacket;                                                                              // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                                    // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                            // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [96:0] addr_router_src_data;                                                                                     // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire  [53:0] addr_router_src_channel;                                                                                  // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                                    // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                             // rsp_xbar_mux:src_endofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                                   // rsp_xbar_mux:src_valid -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                           // rsp_xbar_mux:src_startofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [96:0] rsp_xbar_mux_src_data;                                                                                    // rsp_xbar_mux:src_data -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [53:0] rsp_xbar_mux_src_channel;                                                                                 // rsp_xbar_mux:src_channel -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_src_ready;                                                                                   // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                                          // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                                // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                                        // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [96:0] addr_router_001_src_data;                                                                                 // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire  [53:0] addr_router_001_src_channel;                                                                              // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                                // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                         // rsp_xbar_mux_001:src_endofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                               // rsp_xbar_mux_001:src_valid -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                       // rsp_xbar_mux_001:src_startofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [96:0] rsp_xbar_mux_001_src_data;                                                                                // rsp_xbar_mux_001:src_data -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [53:0] rsp_xbar_mux_001_src_channel;                                                                             // rsp_xbar_mux_001:src_channel -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                               // cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire         addr_router_002_src_endofpacket;                                                                          // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire         addr_router_002_src_valid;                                                                                // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire         addr_router_002_src_startofpacket;                                                                        // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [96:0] addr_router_002_src_data;                                                                                 // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire  [53:0] addr_router_002_src_channel;                                                                              // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire         addr_router_002_src_ready;                                                                                // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire         rsp_xbar_mux_002_src_endofpacket;                                                                         // rsp_xbar_mux_002:src_endofpacket -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_002_src_valid;                                                                               // rsp_xbar_mux_002:src_valid -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_002_src_startofpacket;                                                                       // rsp_xbar_mux_002:src_startofpacket -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [96:0] rsp_xbar_mux_002_src_data;                                                                                // rsp_xbar_mux_002:src_data -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [53:0] rsp_xbar_mux_002_src_channel;                                                                             // rsp_xbar_mux_002:src_channel -> cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_002_src_ready;                                                                               // cpu_1_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_002:src_ready
	wire         addr_router_003_src_endofpacket;                                                                          // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire         addr_router_003_src_valid;                                                                                // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire         addr_router_003_src_startofpacket;                                                                        // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [96:0] addr_router_003_src_data;                                                                                 // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire  [53:0] addr_router_003_src_channel;                                                                              // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire         addr_router_003_src_ready;                                                                                // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire         rsp_xbar_mux_003_src_endofpacket;                                                                         // rsp_xbar_mux_003:src_endofpacket -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_003_src_valid;                                                                               // rsp_xbar_mux_003:src_valid -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_003_src_startofpacket;                                                                       // rsp_xbar_mux_003:src_startofpacket -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [96:0] rsp_xbar_mux_003_src_data;                                                                                // rsp_xbar_mux_003:src_data -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [53:0] rsp_xbar_mux_003_src_channel;                                                                             // rsp_xbar_mux_003:src_channel -> cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_003_src_ready;                                                                               // cpu_1_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_003:src_ready
	wire         addr_router_004_src_endofpacket;                                                                          // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire         addr_router_004_src_valid;                                                                                // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire         addr_router_004_src_startofpacket;                                                                        // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [96:0] addr_router_004_src_data;                                                                                 // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire  [53:0] addr_router_004_src_channel;                                                                              // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire         addr_router_004_src_ready;                                                                                // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire         rsp_xbar_mux_004_src_endofpacket;                                                                         // rsp_xbar_mux_004:src_endofpacket -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_004_src_valid;                                                                               // rsp_xbar_mux_004:src_valid -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_004_src_startofpacket;                                                                       // rsp_xbar_mux_004:src_startofpacket -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [96:0] rsp_xbar_mux_004_src_data;                                                                                // rsp_xbar_mux_004:src_data -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [53:0] rsp_xbar_mux_004_src_channel;                                                                             // rsp_xbar_mux_004:src_channel -> cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_004_src_ready;                                                                               // cpu_2_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_004:src_ready
	wire         addr_router_005_src_endofpacket;                                                                          // addr_router_005:src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire         addr_router_005_src_valid;                                                                                // addr_router_005:src_valid -> cmd_xbar_demux_005:sink_valid
	wire         addr_router_005_src_startofpacket;                                                                        // addr_router_005:src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire  [96:0] addr_router_005_src_data;                                                                                 // addr_router_005:src_data -> cmd_xbar_demux_005:sink_data
	wire  [53:0] addr_router_005_src_channel;                                                                              // addr_router_005:src_channel -> cmd_xbar_demux_005:sink_channel
	wire         addr_router_005_src_ready;                                                                                // cmd_xbar_demux_005:sink_ready -> addr_router_005:src_ready
	wire         rsp_xbar_mux_005_src_endofpacket;                                                                         // rsp_xbar_mux_005:src_endofpacket -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_005_src_valid;                                                                               // rsp_xbar_mux_005:src_valid -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_005_src_startofpacket;                                                                       // rsp_xbar_mux_005:src_startofpacket -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [96:0] rsp_xbar_mux_005_src_data;                                                                                // rsp_xbar_mux_005:src_data -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [53:0] rsp_xbar_mux_005_src_channel;                                                                             // rsp_xbar_mux_005:src_channel -> cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_005_src_ready;                                                                               // cpu_2_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_005:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                             // cmd_xbar_mux:src_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                                   // cmd_xbar_mux:src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                           // cmd_xbar_mux:src_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_src_data;                                                                                    // cmd_xbar_mux:src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_src_channel;                                                                                 // cmd_xbar_mux:src_channel -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                                   // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                                // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                      // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                              // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [96:0] id_router_src_data;                                                                                       // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [53:0] id_router_src_channel;                                                                                    // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                      // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                         // cmd_xbar_mux_001:src_endofpacket -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                               // cmd_xbar_mux_001:src_valid -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                       // cmd_xbar_mux_001:src_startofpacket -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_001_src_data;                                                                                // cmd_xbar_mux_001:src_data -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_001_src_channel;                                                                             // cmd_xbar_mux_001:src_channel -> onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                               // onchip_memory_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                            // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                                  // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                          // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [96:0] id_router_001_src_data;                                                                                   // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire  [53:0] id_router_001_src_channel;                                                                                // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                                  // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                         // cmd_xbar_mux_002:src_endofpacket -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                               // cmd_xbar_mux_002:src_valid -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                       // cmd_xbar_mux_002:src_startofpacket -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_002_src_data;                                                                                // cmd_xbar_mux_002:src_data -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_002_src_channel;                                                                             // cmd_xbar_mux_002:src_channel -> onchip_shared_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                               // onchip_shared_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                            // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                                  // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                          // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [96:0] id_router_002_src_data;                                                                                   // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire  [53:0] id_router_002_src_channel;                                                                                // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                                  // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_001_src3_ready;                                                                            // timer_0_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire         id_router_003_src_endofpacket;                                                                            // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                                  // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                          // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [96:0] id_router_003_src_data;                                                                                   // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire  [53:0] id_router_003_src_channel;                                                                                // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                                  // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_001_src4_ready;                                                                            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire         id_router_004_src_endofpacket;                                                                            // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                                  // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                          // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [96:0] id_router_004_src_data;                                                                                   // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire  [53:0] id_router_004_src_channel;                                                                                // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                                  // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_mux_005_src_endofpacket;                                                                         // cmd_xbar_mux_005:src_endofpacket -> mutex_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_005_src_valid;                                                                               // cmd_xbar_mux_005:src_valid -> mutex_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_005_src_startofpacket;                                                                       // cmd_xbar_mux_005:src_startofpacket -> mutex_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_005_src_data;                                                                                // cmd_xbar_mux_005:src_data -> mutex_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_005_src_channel;                                                                             // cmd_xbar_mux_005:src_channel -> mutex_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_005_src_ready;                                                                               // mutex_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	wire         id_router_005_src_endofpacket;                                                                            // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                                  // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                          // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [96:0] id_router_005_src_data;                                                                                   // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [53:0] id_router_005_src_channel;                                                                                // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                                  // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_mux_006_src_endofpacket;                                                                         // cmd_xbar_mux_006:src_endofpacket -> mutex_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_006_src_valid;                                                                               // cmd_xbar_mux_006:src_valid -> mutex_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_006_src_startofpacket;                                                                       // cmd_xbar_mux_006:src_startofpacket -> mutex_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_006_src_data;                                                                                // cmd_xbar_mux_006:src_data -> mutex_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_006_src_channel;                                                                             // cmd_xbar_mux_006:src_channel -> mutex_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_006_src_ready;                                                                               // mutex_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_006:src_ready
	wire         id_router_006_src_endofpacket;                                                                            // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                                  // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                          // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [96:0] id_router_006_src_data;                                                                                   // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire  [53:0] id_router_006_src_channel;                                                                                // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                                  // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_mux_007_src_endofpacket;                                                                         // cmd_xbar_mux_007:src_endofpacket -> mutex_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_007_src_valid;                                                                               // cmd_xbar_mux_007:src_valid -> mutex_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_007_src_startofpacket;                                                                       // cmd_xbar_mux_007:src_startofpacket -> mutex_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_007_src_data;                                                                                // cmd_xbar_mux_007:src_data -> mutex_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_007_src_channel;                                                                             // cmd_xbar_mux_007:src_channel -> mutex_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_007_src_ready;                                                                               // mutex_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_007:src_ready
	wire         id_router_007_src_endofpacket;                                                                            // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                                  // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                          // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [96:0] id_router_007_src_data;                                                                                   // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire  [53:0] id_router_007_src_channel;                                                                                // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                                  // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_mux_008_src_endofpacket;                                                                         // cmd_xbar_mux_008:src_endofpacket -> mutex_3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_008_src_valid;                                                                               // cmd_xbar_mux_008:src_valid -> mutex_3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_008_src_startofpacket;                                                                       // cmd_xbar_mux_008:src_startofpacket -> mutex_3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_008_src_data;                                                                                // cmd_xbar_mux_008:src_data -> mutex_3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_008_src_channel;                                                                             // cmd_xbar_mux_008:src_channel -> mutex_3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_008_src_ready;                                                                               // mutex_3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_008:src_ready
	wire         id_router_008_src_endofpacket;                                                                            // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                                  // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                          // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [96:0] id_router_008_src_data;                                                                                   // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire  [53:0] id_router_008_src_channel;                                                                                // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                                  // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_mux_009_src_endofpacket;                                                                         // cmd_xbar_mux_009:src_endofpacket -> mutex_4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_009_src_valid;                                                                               // cmd_xbar_mux_009:src_valid -> mutex_4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_009_src_startofpacket;                                                                       // cmd_xbar_mux_009:src_startofpacket -> mutex_4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_009_src_data;                                                                                // cmd_xbar_mux_009:src_data -> mutex_4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_009_src_channel;                                                                             // cmd_xbar_mux_009:src_channel -> mutex_4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_009_src_ready;                                                                               // mutex_4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	wire         id_router_009_src_endofpacket;                                                                            // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         id_router_009_src_valid;                                                                                  // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire         id_router_009_src_startofpacket;                                                                          // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [96:0] id_router_009_src_data;                                                                                   // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire  [53:0] id_router_009_src_channel;                                                                                // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire         id_router_009_src_ready;                                                                                  // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire         cmd_xbar_mux_010_src_endofpacket;                                                                         // cmd_xbar_mux_010:src_endofpacket -> mutex_5_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_010_src_valid;                                                                               // cmd_xbar_mux_010:src_valid -> mutex_5_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_010_src_startofpacket;                                                                       // cmd_xbar_mux_010:src_startofpacket -> mutex_5_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_010_src_data;                                                                                // cmd_xbar_mux_010:src_data -> mutex_5_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_010_src_channel;                                                                             // cmd_xbar_mux_010:src_channel -> mutex_5_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_010_src_ready;                                                                               // mutex_5_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_010:src_ready
	wire         id_router_010_src_endofpacket;                                                                            // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         id_router_010_src_valid;                                                                                  // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire         id_router_010_src_startofpacket;                                                                          // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [96:0] id_router_010_src_data;                                                                                   // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire  [53:0] id_router_010_src_channel;                                                                                // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire         id_router_010_src_ready;                                                                                  // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire         cmd_xbar_demux_001_src11_ready;                                                                           // fifo_0_to_1_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire         id_router_011_src_endofpacket;                                                                            // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire         id_router_011_src_valid;                                                                                  // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire         id_router_011_src_startofpacket;                                                                          // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [96:0] id_router_011_src_data;                                                                                   // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire  [53:0] id_router_011_src_channel;                                                                                // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire         id_router_011_src_ready;                                                                                  // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire         cmd_xbar_demux_001_src12_ready;                                                                           // fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire         id_router_012_src_endofpacket;                                                                            // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire         id_router_012_src_valid;                                                                                  // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire         id_router_012_src_startofpacket;                                                                          // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [96:0] id_router_012_src_data;                                                                                   // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire  [53:0] id_router_012_src_channel;                                                                                // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire         id_router_012_src_ready;                                                                                  // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire         cmd_xbar_demux_001_src13_ready;                                                                           // fifo_0_to_2_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	wire         id_router_013_src_endofpacket;                                                                            // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire         id_router_013_src_valid;                                                                                  // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire         id_router_013_src_startofpacket;                                                                          // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [96:0] id_router_013_src_data;                                                                                   // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire  [53:0] id_router_013_src_channel;                                                                                // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire         id_router_013_src_ready;                                                                                  // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire         cmd_xbar_demux_001_src14_ready;                                                                           // fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	wire         id_router_014_src_endofpacket;                                                                            // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire         id_router_014_src_valid;                                                                                  // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire         id_router_014_src_startofpacket;                                                                          // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [96:0] id_router_014_src_data;                                                                                   // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire  [53:0] id_router_014_src_channel;                                                                                // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire         id_router_014_src_ready;                                                                                  // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire         cmd_xbar_demux_001_src15_ready;                                                                           // fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	wire         id_router_015_src_endofpacket;                                                                            // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire         id_router_015_src_valid;                                                                                  // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire         id_router_015_src_startofpacket;                                                                          // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [96:0] id_router_015_src_data;                                                                                   // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire  [53:0] id_router_015_src_channel;                                                                                // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire         id_router_015_src_ready;                                                                                  // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire         cmd_xbar_demux_001_src16_ready;                                                                           // fifo_1_to_0_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src16_ready
	wire         id_router_016_src_endofpacket;                                                                            // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire         id_router_016_src_valid;                                                                                  // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire         id_router_016_src_startofpacket;                                                                          // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [96:0] id_router_016_src_data;                                                                                   // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire  [53:0] id_router_016_src_channel;                                                                                // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire         id_router_016_src_ready;                                                                                  // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire         cmd_xbar_demux_001_src17_ready;                                                                           // fifo_2_to_0_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src17_ready
	wire         id_router_017_src_endofpacket;                                                                            // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire         id_router_017_src_valid;                                                                                  // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire         id_router_017_src_startofpacket;                                                                          // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [96:0] id_router_017_src_data;                                                                                   // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire  [53:0] id_router_017_src_channel;                                                                                // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire         id_router_017_src_ready;                                                                                  // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire         cmd_xbar_demux_001_src18_ready;                                                                           // fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src18_ready
	wire         id_router_018_src_endofpacket;                                                                            // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire         id_router_018_src_valid;                                                                                  // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire         id_router_018_src_startofpacket;                                                                          // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [96:0] id_router_018_src_data;                                                                                   // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire  [53:0] id_router_018_src_channel;                                                                                // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire         id_router_018_src_ready;                                                                                  // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire         cmd_xbar_mux_019_src_endofpacket;                                                                         // cmd_xbar_mux_019:src_endofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_019_src_valid;                                                                               // cmd_xbar_mux_019:src_valid -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_019_src_startofpacket;                                                                       // cmd_xbar_mux_019:src_startofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_019_src_data;                                                                                // cmd_xbar_mux_019:src_data -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_019_src_channel;                                                                             // cmd_xbar_mux_019:src_channel -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_019_src_ready;                                                                               // red_leds_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_019:src_ready
	wire         id_router_019_src_endofpacket;                                                                            // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire         id_router_019_src_valid;                                                                                  // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire         id_router_019_src_startofpacket;                                                                          // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [96:0] id_router_019_src_data;                                                                                   // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire  [53:0] id_router_019_src_channel;                                                                                // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire         id_router_019_src_ready;                                                                                  // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire         cmd_xbar_mux_020_src_endofpacket;                                                                         // cmd_xbar_mux_020:src_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_020_src_valid;                                                                               // cmd_xbar_mux_020:src_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_020_src_startofpacket;                                                                       // cmd_xbar_mux_020:src_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_020_src_data;                                                                                // cmd_xbar_mux_020:src_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_020_src_channel;                                                                             // cmd_xbar_mux_020:src_channel -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_020_src_ready;                                                                               // green_leds_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_020:src_ready
	wire         id_router_020_src_endofpacket;                                                                            // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire         id_router_020_src_valid;                                                                                  // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire         id_router_020_src_startofpacket;                                                                          // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [96:0] id_router_020_src_data;                                                                                   // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire  [53:0] id_router_020_src_channel;                                                                                // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire         id_router_020_src_ready;                                                                                  // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire         cmd_xbar_mux_021_src_endofpacket;                                                                         // cmd_xbar_mux_021:src_endofpacket -> switches_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_021_src_valid;                                                                               // cmd_xbar_mux_021:src_valid -> switches_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_021_src_startofpacket;                                                                       // cmd_xbar_mux_021:src_startofpacket -> switches_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_021_src_data;                                                                                // cmd_xbar_mux_021:src_data -> switches_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_021_src_channel;                                                                             // cmd_xbar_mux_021:src_channel -> switches_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_021_src_ready;                                                                               // switches_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_021:src_ready
	wire         id_router_021_src_endofpacket;                                                                            // id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire         id_router_021_src_valid;                                                                                  // id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	wire         id_router_021_src_startofpacket;                                                                          // id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [96:0] id_router_021_src_data;                                                                                   // id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	wire  [53:0] id_router_021_src_channel;                                                                                // id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	wire         id_router_021_src_ready;                                                                                  // rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	wire         cmd_xbar_mux_022_src_endofpacket;                                                                         // cmd_xbar_mux_022:src_endofpacket -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_022_src_valid;                                                                               // cmd_xbar_mux_022:src_valid -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_022_src_startofpacket;                                                                       // cmd_xbar_mux_022:src_startofpacket -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_022_src_data;                                                                                // cmd_xbar_mux_022:src_data -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_022_src_channel;                                                                             // cmd_xbar_mux_022:src_channel -> timer_shared_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_022_src_ready;                                                                               // timer_shared_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_022:src_ready
	wire         id_router_022_src_endofpacket;                                                                            // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire         id_router_022_src_valid;                                                                                  // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire         id_router_022_src_startofpacket;                                                                          // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire  [96:0] id_router_022_src_data;                                                                                   // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire  [53:0] id_router_022_src_channel;                                                                                // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire         id_router_022_src_ready;                                                                                  // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire         cmd_xbar_demux_001_src23_ready;                                                                           // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src23_ready
	wire         id_router_023_src_endofpacket;                                                                            // id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire         id_router_023_src_valid;                                                                                  // id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	wire         id_router_023_src_startofpacket;                                                                          // id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire  [96:0] id_router_023_src_data;                                                                                   // id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	wire  [53:0] id_router_023_src_channel;                                                                                // id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	wire         id_router_023_src_ready;                                                                                  // rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	wire         cmd_xbar_demux_001_src24_ready;                                                                           // timer_0_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src24_ready
	wire         id_router_024_src_endofpacket;                                                                            // id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire         id_router_024_src_valid;                                                                                  // id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	wire         id_router_024_src_startofpacket;                                                                          // id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire  [96:0] id_router_024_src_data;                                                                                   // id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	wire  [53:0] id_router_024_src_channel;                                                                                // id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	wire         id_router_024_src_ready;                                                                                  // rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	wire         cmd_xbar_mux_025_src_endofpacket;                                                                         // cmd_xbar_mux_025:src_endofpacket -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_025_src_valid;                                                                               // cmd_xbar_mux_025:src_valid -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_025_src_startofpacket;                                                                       // cmd_xbar_mux_025:src_startofpacket -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_025_src_data;                                                                                // cmd_xbar_mux_025:src_data -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_025_src_channel;                                                                             // cmd_xbar_mux_025:src_channel -> timer_shared_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_025_src_ready;                                                                               // timer_shared_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_025:src_ready
	wire         id_router_025_src_endofpacket;                                                                            // id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	wire         id_router_025_src_valid;                                                                                  // id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	wire         id_router_025_src_startofpacket;                                                                          // id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	wire  [96:0] id_router_025_src_data;                                                                                   // id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	wire  [53:0] id_router_025_src_channel;                                                                                // id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	wire         id_router_025_src_ready;                                                                                  // rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	wire         cmd_xbar_mux_026_src_endofpacket;                                                                         // cmd_xbar_mux_026:src_endofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_026_src_valid;                                                                               // cmd_xbar_mux_026:src_valid -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_026_src_startofpacket;                                                                       // cmd_xbar_mux_026:src_startofpacket -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_026_src_data;                                                                                // cmd_xbar_mux_026:src_data -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_026_src_channel;                                                                             // cmd_xbar_mux_026:src_channel -> cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_026_src_ready;                                                                               // cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_026:src_ready
	wire         id_router_026_src_endofpacket;                                                                            // id_router_026:src_endofpacket -> rsp_xbar_demux_026:sink_endofpacket
	wire         id_router_026_src_valid;                                                                                  // id_router_026:src_valid -> rsp_xbar_demux_026:sink_valid
	wire         id_router_026_src_startofpacket;                                                                          // id_router_026:src_startofpacket -> rsp_xbar_demux_026:sink_startofpacket
	wire  [96:0] id_router_026_src_data;                                                                                   // id_router_026:src_data -> rsp_xbar_demux_026:sink_data
	wire  [53:0] id_router_026_src_channel;                                                                                // id_router_026:src_channel -> rsp_xbar_demux_026:sink_channel
	wire         id_router_026_src_ready;                                                                                  // rsp_xbar_demux_026:sink_ready -> id_router_026:src_ready
	wire         cmd_xbar_mux_027_src_endofpacket;                                                                         // cmd_xbar_mux_027:src_endofpacket -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_027_src_valid;                                                                               // cmd_xbar_mux_027:src_valid -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_027_src_startofpacket;                                                                       // cmd_xbar_mux_027:src_startofpacket -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_027_src_data;                                                                                // cmd_xbar_mux_027:src_data -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_027_src_channel;                                                                             // cmd_xbar_mux_027:src_channel -> onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_027_src_ready;                                                                               // onchip_memory_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_027:src_ready
	wire         id_router_027_src_endofpacket;                                                                            // id_router_027:src_endofpacket -> rsp_xbar_demux_027:sink_endofpacket
	wire         id_router_027_src_valid;                                                                                  // id_router_027:src_valid -> rsp_xbar_demux_027:sink_valid
	wire         id_router_027_src_startofpacket;                                                                          // id_router_027:src_startofpacket -> rsp_xbar_demux_027:sink_startofpacket
	wire  [96:0] id_router_027_src_data;                                                                                   // id_router_027:src_data -> rsp_xbar_demux_027:sink_data
	wire  [53:0] id_router_027_src_channel;                                                                                // id_router_027:src_channel -> rsp_xbar_demux_027:sink_channel
	wire         id_router_027_src_ready;                                                                                  // rsp_xbar_demux_027:sink_ready -> id_router_027:src_ready
	wire         cmd_xbar_demux_002_src14_ready;                                                                           // timer_1_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src14_ready
	wire         id_router_028_src_endofpacket;                                                                            // id_router_028:src_endofpacket -> rsp_xbar_demux_028:sink_endofpacket
	wire         id_router_028_src_valid;                                                                                  // id_router_028:src_valid -> rsp_xbar_demux_028:sink_valid
	wire         id_router_028_src_startofpacket;                                                                          // id_router_028:src_startofpacket -> rsp_xbar_demux_028:sink_startofpacket
	wire  [96:0] id_router_028_src_data;                                                                                   // id_router_028:src_data -> rsp_xbar_demux_028:sink_data
	wire  [53:0] id_router_028_src_channel;                                                                                // id_router_028:src_channel -> rsp_xbar_demux_028:sink_channel
	wire         id_router_028_src_ready;                                                                                  // rsp_xbar_demux_028:sink_ready -> id_router_028:src_ready
	wire         cmd_xbar_demux_002_src15_ready;                                                                           // jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src15_ready
	wire         id_router_029_src_endofpacket;                                                                            // id_router_029:src_endofpacket -> rsp_xbar_demux_029:sink_endofpacket
	wire         id_router_029_src_valid;                                                                                  // id_router_029:src_valid -> rsp_xbar_demux_029:sink_valid
	wire         id_router_029_src_startofpacket;                                                                          // id_router_029:src_startofpacket -> rsp_xbar_demux_029:sink_startofpacket
	wire  [96:0] id_router_029_src_data;                                                                                   // id_router_029:src_data -> rsp_xbar_demux_029:sink_data
	wire  [53:0] id_router_029_src_channel;                                                                                // id_router_029:src_channel -> rsp_xbar_demux_029:sink_channel
	wire         id_router_029_src_ready;                                                                                  // rsp_xbar_demux_029:sink_ready -> id_router_029:src_ready
	wire         cmd_xbar_demux_002_src16_ready;                                                                           // fifo_0_to_1_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src16_ready
	wire         id_router_030_src_endofpacket;                                                                            // id_router_030:src_endofpacket -> rsp_xbar_demux_030:sink_endofpacket
	wire         id_router_030_src_valid;                                                                                  // id_router_030:src_valid -> rsp_xbar_demux_030:sink_valid
	wire         id_router_030_src_startofpacket;                                                                          // id_router_030:src_startofpacket -> rsp_xbar_demux_030:sink_startofpacket
	wire  [96:0] id_router_030_src_data;                                                                                   // id_router_030:src_data -> rsp_xbar_demux_030:sink_data
	wire  [53:0] id_router_030_src_channel;                                                                                // id_router_030:src_channel -> rsp_xbar_demux_030:sink_channel
	wire         id_router_030_src_ready;                                                                                  // rsp_xbar_demux_030:sink_ready -> id_router_030:src_ready
	wire         cmd_xbar_demux_002_src17_ready;                                                                           // fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src17_ready
	wire         id_router_031_src_endofpacket;                                                                            // id_router_031:src_endofpacket -> rsp_xbar_demux_031:sink_endofpacket
	wire         id_router_031_src_valid;                                                                                  // id_router_031:src_valid -> rsp_xbar_demux_031:sink_valid
	wire         id_router_031_src_startofpacket;                                                                          // id_router_031:src_startofpacket -> rsp_xbar_demux_031:sink_startofpacket
	wire  [96:0] id_router_031_src_data;                                                                                   // id_router_031:src_data -> rsp_xbar_demux_031:sink_data
	wire  [53:0] id_router_031_src_channel;                                                                                // id_router_031:src_channel -> rsp_xbar_demux_031:sink_channel
	wire         id_router_031_src_ready;                                                                                  // rsp_xbar_demux_031:sink_ready -> id_router_031:src_ready
	wire         cmd_xbar_demux_002_src18_ready;                                                                           // fifo_1_to_0_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src18_ready
	wire         id_router_032_src_endofpacket;                                                                            // id_router_032:src_endofpacket -> rsp_xbar_demux_032:sink_endofpacket
	wire         id_router_032_src_valid;                                                                                  // id_router_032:src_valid -> rsp_xbar_demux_032:sink_valid
	wire         id_router_032_src_startofpacket;                                                                          // id_router_032:src_startofpacket -> rsp_xbar_demux_032:sink_startofpacket
	wire  [96:0] id_router_032_src_data;                                                                                   // id_router_032:src_data -> rsp_xbar_demux_032:sink_data
	wire  [53:0] id_router_032_src_channel;                                                                                // id_router_032:src_channel -> rsp_xbar_demux_032:sink_channel
	wire         id_router_032_src_ready;                                                                                  // rsp_xbar_demux_032:sink_ready -> id_router_032:src_ready
	wire         cmd_xbar_demux_002_src19_ready;                                                                           // fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src19_ready
	wire         id_router_033_src_endofpacket;                                                                            // id_router_033:src_endofpacket -> rsp_xbar_demux_033:sink_endofpacket
	wire         id_router_033_src_valid;                                                                                  // id_router_033:src_valid -> rsp_xbar_demux_033:sink_valid
	wire         id_router_033_src_startofpacket;                                                                          // id_router_033:src_startofpacket -> rsp_xbar_demux_033:sink_startofpacket
	wire  [96:0] id_router_033_src_data;                                                                                   // id_router_033:src_data -> rsp_xbar_demux_033:sink_data
	wire  [53:0] id_router_033_src_channel;                                                                                // id_router_033:src_channel -> rsp_xbar_demux_033:sink_channel
	wire         id_router_033_src_ready;                                                                                  // rsp_xbar_demux_033:sink_ready -> id_router_033:src_ready
	wire         cmd_xbar_demux_002_src20_ready;                                                                           // fifo_1_to_2_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src20_ready
	wire         id_router_034_src_endofpacket;                                                                            // id_router_034:src_endofpacket -> rsp_xbar_demux_034:sink_endofpacket
	wire         id_router_034_src_valid;                                                                                  // id_router_034:src_valid -> rsp_xbar_demux_034:sink_valid
	wire         id_router_034_src_startofpacket;                                                                          // id_router_034:src_startofpacket -> rsp_xbar_demux_034:sink_startofpacket
	wire  [96:0] id_router_034_src_data;                                                                                   // id_router_034:src_data -> rsp_xbar_demux_034:sink_data
	wire  [53:0] id_router_034_src_channel;                                                                                // id_router_034:src_channel -> rsp_xbar_demux_034:sink_channel
	wire         id_router_034_src_ready;                                                                                  // rsp_xbar_demux_034:sink_ready -> id_router_034:src_ready
	wire         cmd_xbar_demux_002_src21_ready;                                                                           // fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src21_ready
	wire         id_router_035_src_endofpacket;                                                                            // id_router_035:src_endofpacket -> rsp_xbar_demux_035:sink_endofpacket
	wire         id_router_035_src_valid;                                                                                  // id_router_035:src_valid -> rsp_xbar_demux_035:sink_valid
	wire         id_router_035_src_startofpacket;                                                                          // id_router_035:src_startofpacket -> rsp_xbar_demux_035:sink_startofpacket
	wire  [96:0] id_router_035_src_data;                                                                                   // id_router_035:src_data -> rsp_xbar_demux_035:sink_data
	wire  [53:0] id_router_035_src_channel;                                                                                // id_router_035:src_channel -> rsp_xbar_demux_035:sink_channel
	wire         id_router_035_src_ready;                                                                                  // rsp_xbar_demux_035:sink_ready -> id_router_035:src_ready
	wire         cmd_xbar_demux_002_src22_ready;                                                                           // fifo_2_to_1_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src22_ready
	wire         id_router_036_src_endofpacket;                                                                            // id_router_036:src_endofpacket -> rsp_xbar_demux_036:sink_endofpacket
	wire         id_router_036_src_valid;                                                                                  // id_router_036:src_valid -> rsp_xbar_demux_036:sink_valid
	wire         id_router_036_src_startofpacket;                                                                          // id_router_036:src_startofpacket -> rsp_xbar_demux_036:sink_startofpacket
	wire  [96:0] id_router_036_src_data;                                                                                   // id_router_036:src_data -> rsp_xbar_demux_036:sink_data
	wire  [53:0] id_router_036_src_channel;                                                                                // id_router_036:src_channel -> rsp_xbar_demux_036:sink_channel
	wire         id_router_036_src_ready;                                                                                  // rsp_xbar_demux_036:sink_ready -> id_router_036:src_ready
	wire         cmd_xbar_demux_002_src23_ready;                                                                           // fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src23_ready
	wire         id_router_037_src_endofpacket;                                                                            // id_router_037:src_endofpacket -> rsp_xbar_demux_037:sink_endofpacket
	wire         id_router_037_src_valid;                                                                                  // id_router_037:src_valid -> rsp_xbar_demux_037:sink_valid
	wire         id_router_037_src_startofpacket;                                                                          // id_router_037:src_startofpacket -> rsp_xbar_demux_037:sink_startofpacket
	wire  [96:0] id_router_037_src_data;                                                                                   // id_router_037:src_data -> rsp_xbar_demux_037:sink_data
	wire  [53:0] id_router_037_src_channel;                                                                                // id_router_037:src_channel -> rsp_xbar_demux_037:sink_channel
	wire         id_router_037_src_ready;                                                                                  // rsp_xbar_demux_037:sink_ready -> id_router_037:src_ready
	wire         cmd_xbar_demux_002_src24_ready;                                                                           // performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src24_ready
	wire         id_router_038_src_endofpacket;                                                                            // id_router_038:src_endofpacket -> rsp_xbar_demux_038:sink_endofpacket
	wire         id_router_038_src_valid;                                                                                  // id_router_038:src_valid -> rsp_xbar_demux_038:sink_valid
	wire         id_router_038_src_startofpacket;                                                                          // id_router_038:src_startofpacket -> rsp_xbar_demux_038:sink_startofpacket
	wire  [96:0] id_router_038_src_data;                                                                                   // id_router_038:src_data -> rsp_xbar_demux_038:sink_data
	wire  [53:0] id_router_038_src_channel;                                                                                // id_router_038:src_channel -> rsp_xbar_demux_038:sink_channel
	wire         id_router_038_src_ready;                                                                                  // rsp_xbar_demux_038:sink_ready -> id_router_038:src_ready
	wire         cmd_xbar_demux_002_src25_ready;                                                                           // timer_1_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src25_ready
	wire         id_router_039_src_endofpacket;                                                                            // id_router_039:src_endofpacket -> rsp_xbar_demux_039:sink_endofpacket
	wire         id_router_039_src_valid;                                                                                  // id_router_039:src_valid -> rsp_xbar_demux_039:sink_valid
	wire         id_router_039_src_startofpacket;                                                                          // id_router_039:src_startofpacket -> rsp_xbar_demux_039:sink_startofpacket
	wire  [96:0] id_router_039_src_data;                                                                                   // id_router_039:src_data -> rsp_xbar_demux_039:sink_data
	wire  [53:0] id_router_039_src_channel;                                                                                // id_router_039:src_channel -> rsp_xbar_demux_039:sink_channel
	wire         id_router_039_src_ready;                                                                                  // rsp_xbar_demux_039:sink_ready -> id_router_039:src_ready
	wire         cmd_xbar_mux_040_src_endofpacket;                                                                         // cmd_xbar_mux_040:src_endofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_040_src_valid;                                                                               // cmd_xbar_mux_040:src_valid -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_040_src_startofpacket;                                                                       // cmd_xbar_mux_040:src_startofpacket -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_040_src_data;                                                                                // cmd_xbar_mux_040:src_data -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_040_src_channel;                                                                             // cmd_xbar_mux_040:src_channel -> cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_040_src_ready;                                                                               // cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_040:src_ready
	wire         id_router_040_src_endofpacket;                                                                            // id_router_040:src_endofpacket -> rsp_xbar_demux_040:sink_endofpacket
	wire         id_router_040_src_valid;                                                                                  // id_router_040:src_valid -> rsp_xbar_demux_040:sink_valid
	wire         id_router_040_src_startofpacket;                                                                          // id_router_040:src_startofpacket -> rsp_xbar_demux_040:sink_startofpacket
	wire  [96:0] id_router_040_src_data;                                                                                   // id_router_040:src_data -> rsp_xbar_demux_040:sink_data
	wire  [53:0] id_router_040_src_channel;                                                                                // id_router_040:src_channel -> rsp_xbar_demux_040:sink_channel
	wire         id_router_040_src_ready;                                                                                  // rsp_xbar_demux_040:sink_ready -> id_router_040:src_ready
	wire         cmd_xbar_mux_041_src_endofpacket;                                                                         // cmd_xbar_mux_041:src_endofpacket -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_041_src_valid;                                                                               // cmd_xbar_mux_041:src_valid -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_041_src_startofpacket;                                                                       // cmd_xbar_mux_041:src_startofpacket -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [96:0] cmd_xbar_mux_041_src_data;                                                                                // cmd_xbar_mux_041:src_data -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [53:0] cmd_xbar_mux_041_src_channel;                                                                             // cmd_xbar_mux_041:src_channel -> onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_041_src_ready;                                                                               // onchip_memory_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_041:src_ready
	wire         id_router_041_src_endofpacket;                                                                            // id_router_041:src_endofpacket -> rsp_xbar_demux_041:sink_endofpacket
	wire         id_router_041_src_valid;                                                                                  // id_router_041:src_valid -> rsp_xbar_demux_041:sink_valid
	wire         id_router_041_src_startofpacket;                                                                          // id_router_041:src_startofpacket -> rsp_xbar_demux_041:sink_startofpacket
	wire  [96:0] id_router_041_src_data;                                                                                   // id_router_041:src_data -> rsp_xbar_demux_041:sink_data
	wire  [53:0] id_router_041_src_channel;                                                                                // id_router_041:src_channel -> rsp_xbar_demux_041:sink_channel
	wire         id_router_041_src_ready;                                                                                  // rsp_xbar_demux_041:sink_ready -> id_router_041:src_ready
	wire         cmd_xbar_demux_004_src14_ready;                                                                           // timer_2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src14_ready
	wire         id_router_042_src_endofpacket;                                                                            // id_router_042:src_endofpacket -> rsp_xbar_demux_042:sink_endofpacket
	wire         id_router_042_src_valid;                                                                                  // id_router_042:src_valid -> rsp_xbar_demux_042:sink_valid
	wire         id_router_042_src_startofpacket;                                                                          // id_router_042:src_startofpacket -> rsp_xbar_demux_042:sink_startofpacket
	wire  [96:0] id_router_042_src_data;                                                                                   // id_router_042:src_data -> rsp_xbar_demux_042:sink_data
	wire  [53:0] id_router_042_src_channel;                                                                                // id_router_042:src_channel -> rsp_xbar_demux_042:sink_channel
	wire         id_router_042_src_ready;                                                                                  // rsp_xbar_demux_042:sink_ready -> id_router_042:src_ready
	wire         cmd_xbar_demux_004_src15_ready;                                                                           // jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src15_ready
	wire         id_router_043_src_endofpacket;                                                                            // id_router_043:src_endofpacket -> rsp_xbar_demux_043:sink_endofpacket
	wire         id_router_043_src_valid;                                                                                  // id_router_043:src_valid -> rsp_xbar_demux_043:sink_valid
	wire         id_router_043_src_startofpacket;                                                                          // id_router_043:src_startofpacket -> rsp_xbar_demux_043:sink_startofpacket
	wire  [96:0] id_router_043_src_data;                                                                                   // id_router_043:src_data -> rsp_xbar_demux_043:sink_data
	wire  [53:0] id_router_043_src_channel;                                                                                // id_router_043:src_channel -> rsp_xbar_demux_043:sink_channel
	wire         id_router_043_src_ready;                                                                                  // rsp_xbar_demux_043:sink_ready -> id_router_043:src_ready
	wire         cmd_xbar_demux_004_src16_ready;                                                                           // fifo_0_to_2_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src16_ready
	wire         id_router_044_src_endofpacket;                                                                            // id_router_044:src_endofpacket -> rsp_xbar_demux_044:sink_endofpacket
	wire         id_router_044_src_valid;                                                                                  // id_router_044:src_valid -> rsp_xbar_demux_044:sink_valid
	wire         id_router_044_src_startofpacket;                                                                          // id_router_044:src_startofpacket -> rsp_xbar_demux_044:sink_startofpacket
	wire  [96:0] id_router_044_src_data;                                                                                   // id_router_044:src_data -> rsp_xbar_demux_044:sink_data
	wire  [53:0] id_router_044_src_channel;                                                                                // id_router_044:src_channel -> rsp_xbar_demux_044:sink_channel
	wire         id_router_044_src_ready;                                                                                  // rsp_xbar_demux_044:sink_ready -> id_router_044:src_ready
	wire         cmd_xbar_demux_004_src17_ready;                                                                           // fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src17_ready
	wire         id_router_045_src_endofpacket;                                                                            // id_router_045:src_endofpacket -> rsp_xbar_demux_045:sink_endofpacket
	wire         id_router_045_src_valid;                                                                                  // id_router_045:src_valid -> rsp_xbar_demux_045:sink_valid
	wire         id_router_045_src_startofpacket;                                                                          // id_router_045:src_startofpacket -> rsp_xbar_demux_045:sink_startofpacket
	wire  [96:0] id_router_045_src_data;                                                                                   // id_router_045:src_data -> rsp_xbar_demux_045:sink_data
	wire  [53:0] id_router_045_src_channel;                                                                                // id_router_045:src_channel -> rsp_xbar_demux_045:sink_channel
	wire         id_router_045_src_ready;                                                                                  // rsp_xbar_demux_045:sink_ready -> id_router_045:src_ready
	wire         cmd_xbar_demux_004_src18_ready;                                                                           // fifo_1_to_2_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src18_ready
	wire         id_router_046_src_endofpacket;                                                                            // id_router_046:src_endofpacket -> rsp_xbar_demux_046:sink_endofpacket
	wire         id_router_046_src_valid;                                                                                  // id_router_046:src_valid -> rsp_xbar_demux_046:sink_valid
	wire         id_router_046_src_startofpacket;                                                                          // id_router_046:src_startofpacket -> rsp_xbar_demux_046:sink_startofpacket
	wire  [96:0] id_router_046_src_data;                                                                                   // id_router_046:src_data -> rsp_xbar_demux_046:sink_data
	wire  [53:0] id_router_046_src_channel;                                                                                // id_router_046:src_channel -> rsp_xbar_demux_046:sink_channel
	wire         id_router_046_src_ready;                                                                                  // rsp_xbar_demux_046:sink_ready -> id_router_046:src_ready
	wire         cmd_xbar_demux_004_src19_ready;                                                                           // fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src19_ready
	wire         id_router_047_src_endofpacket;                                                                            // id_router_047:src_endofpacket -> rsp_xbar_demux_047:sink_endofpacket
	wire         id_router_047_src_valid;                                                                                  // id_router_047:src_valid -> rsp_xbar_demux_047:sink_valid
	wire         id_router_047_src_startofpacket;                                                                          // id_router_047:src_startofpacket -> rsp_xbar_demux_047:sink_startofpacket
	wire  [96:0] id_router_047_src_data;                                                                                   // id_router_047:src_data -> rsp_xbar_demux_047:sink_data
	wire  [53:0] id_router_047_src_channel;                                                                                // id_router_047:src_channel -> rsp_xbar_demux_047:sink_channel
	wire         id_router_047_src_ready;                                                                                  // rsp_xbar_demux_047:sink_ready -> id_router_047:src_ready
	wire         cmd_xbar_demux_004_src20_ready;                                                                           // fifo_2_to_0_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src20_ready
	wire         id_router_048_src_endofpacket;                                                                            // id_router_048:src_endofpacket -> rsp_xbar_demux_048:sink_endofpacket
	wire         id_router_048_src_valid;                                                                                  // id_router_048:src_valid -> rsp_xbar_demux_048:sink_valid
	wire         id_router_048_src_startofpacket;                                                                          // id_router_048:src_startofpacket -> rsp_xbar_demux_048:sink_startofpacket
	wire  [96:0] id_router_048_src_data;                                                                                   // id_router_048:src_data -> rsp_xbar_demux_048:sink_data
	wire  [53:0] id_router_048_src_channel;                                                                                // id_router_048:src_channel -> rsp_xbar_demux_048:sink_channel
	wire         id_router_048_src_ready;                                                                                  // rsp_xbar_demux_048:sink_ready -> id_router_048:src_ready
	wire         cmd_xbar_demux_004_src21_ready;                                                                           // fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src21_ready
	wire         id_router_049_src_endofpacket;                                                                            // id_router_049:src_endofpacket -> rsp_xbar_demux_049:sink_endofpacket
	wire         id_router_049_src_valid;                                                                                  // id_router_049:src_valid -> rsp_xbar_demux_049:sink_valid
	wire         id_router_049_src_startofpacket;                                                                          // id_router_049:src_startofpacket -> rsp_xbar_demux_049:sink_startofpacket
	wire  [96:0] id_router_049_src_data;                                                                                   // id_router_049:src_data -> rsp_xbar_demux_049:sink_data
	wire  [53:0] id_router_049_src_channel;                                                                                // id_router_049:src_channel -> rsp_xbar_demux_049:sink_channel
	wire         id_router_049_src_ready;                                                                                  // rsp_xbar_demux_049:sink_ready -> id_router_049:src_ready
	wire         cmd_xbar_demux_004_src22_ready;                                                                           // fifo_2_to_1_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src22_ready
	wire         id_router_050_src_endofpacket;                                                                            // id_router_050:src_endofpacket -> rsp_xbar_demux_050:sink_endofpacket
	wire         id_router_050_src_valid;                                                                                  // id_router_050:src_valid -> rsp_xbar_demux_050:sink_valid
	wire         id_router_050_src_startofpacket;                                                                          // id_router_050:src_startofpacket -> rsp_xbar_demux_050:sink_startofpacket
	wire  [96:0] id_router_050_src_data;                                                                                   // id_router_050:src_data -> rsp_xbar_demux_050:sink_data
	wire  [53:0] id_router_050_src_channel;                                                                                // id_router_050:src_channel -> rsp_xbar_demux_050:sink_channel
	wire         id_router_050_src_ready;                                                                                  // rsp_xbar_demux_050:sink_ready -> id_router_050:src_ready
	wire         cmd_xbar_demux_004_src23_ready;                                                                           // fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src23_ready
	wire         id_router_051_src_endofpacket;                                                                            // id_router_051:src_endofpacket -> rsp_xbar_demux_051:sink_endofpacket
	wire         id_router_051_src_valid;                                                                                  // id_router_051:src_valid -> rsp_xbar_demux_051:sink_valid
	wire         id_router_051_src_startofpacket;                                                                          // id_router_051:src_startofpacket -> rsp_xbar_demux_051:sink_startofpacket
	wire  [96:0] id_router_051_src_data;                                                                                   // id_router_051:src_data -> rsp_xbar_demux_051:sink_data
	wire  [53:0] id_router_051_src_channel;                                                                                // id_router_051:src_channel -> rsp_xbar_demux_051:sink_channel
	wire         id_router_051_src_ready;                                                                                  // rsp_xbar_demux_051:sink_ready -> id_router_051:src_ready
	wire         cmd_xbar_demux_004_src24_ready;                                                                           // performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src24_ready
	wire         id_router_052_src_endofpacket;                                                                            // id_router_052:src_endofpacket -> rsp_xbar_demux_052:sink_endofpacket
	wire         id_router_052_src_valid;                                                                                  // id_router_052:src_valid -> rsp_xbar_demux_052:sink_valid
	wire         id_router_052_src_startofpacket;                                                                          // id_router_052:src_startofpacket -> rsp_xbar_demux_052:sink_startofpacket
	wire  [96:0] id_router_052_src_data;                                                                                   // id_router_052:src_data -> rsp_xbar_demux_052:sink_data
	wire  [53:0] id_router_052_src_channel;                                                                                // id_router_052:src_channel -> rsp_xbar_demux_052:sink_channel
	wire         id_router_052_src_ready;                                                                                  // rsp_xbar_demux_052:sink_ready -> id_router_052:src_ready
	wire         cmd_xbar_demux_004_src25_ready;                                                                           // timer_2_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src25_ready
	wire         id_router_053_src_endofpacket;                                                                            // id_router_053:src_endofpacket -> rsp_xbar_demux_053:sink_endofpacket
	wire         id_router_053_src_valid;                                                                                  // id_router_053:src_valid -> rsp_xbar_demux_053:sink_valid
	wire         id_router_053_src_startofpacket;                                                                          // id_router_053:src_startofpacket -> rsp_xbar_demux_053:sink_startofpacket
	wire  [96:0] id_router_053_src_data;                                                                                   // id_router_053:src_data -> rsp_xbar_demux_053:sink_data
	wire  [53:0] id_router_053_src_channel;                                                                                // id_router_053:src_channel -> rsp_xbar_demux_053:sink_channel
	wire         id_router_053_src_ready;                                                                                  // rsp_xbar_demux_053:sink_ready -> id_router_053:src_ready
	wire         irq_mapper_receiver0_irq;                                                                                 // timer_0_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                                 // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver3_irq;                                                                                 // timer_0_1:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_0_d_irq_irq;                                                                                          // irq_mapper:sender_irq -> cpu_0:d_irq
	wire         irq_mapper_001_receiver0_irq;                                                                             // timer_1_0:irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                                                                             // jtag_uart_1:av_irq -> irq_mapper_001:receiver1_irq
	wire         irq_mapper_001_receiver3_irq;                                                                             // timer_1_1:irq -> irq_mapper_001:receiver3_irq
	wire  [31:0] cpu_1_d_irq_irq;                                                                                          // irq_mapper_001:sender_irq -> cpu_1:d_irq
	wire         irq_mapper_002_receiver0_irq;                                                                             // timer_2_0:irq -> irq_mapper_002:receiver0_irq
	wire         irq_mapper_002_receiver1_irq;                                                                             // jtag_uart_2:av_irq -> irq_mapper_002:receiver1_irq
	wire         irq_mapper_002_receiver3_irq;                                                                             // timer_2_1:irq -> irq_mapper_002:receiver3_irq
	wire  [31:0] cpu_2_d_irq_irq;                                                                                          // irq_mapper_002:sender_irq -> cpu_2:d_irq
	wire         irq_mapper_receiver2_irq;                                                                                 // timer_shared_0:irq -> [irq_mapper:receiver2_irq, irq_mapper_001:receiver2_irq, irq_mapper_002:receiver2_irq]
	wire         irq_mapper_receiver4_irq;                                                                                 // timer_shared_1:irq -> [irq_mapper:receiver4_irq, irq_mapper_001:receiver4_irq, irq_mapper_002:receiver4_irq]

	Core3_cpu_0 cpu_0 (
		.clk                                   (clk_clk),                                                            //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                    //                   reset_n.reset_n
		.d_address                             (cpu_0_data_master_address),                                          //               data_master.address
		.d_byteenable                          (cpu_0_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (cpu_0_data_master_read),                                             //                          .read
		.d_readdata                            (cpu_0_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (cpu_0_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (cpu_0_data_master_write),                                            //                          .write
		.d_writedata                           (cpu_0_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_0_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (cpu_0_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (cpu_0_instruction_master_read),                                      //                          .read
		.i_readdata                            (cpu_0_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (cpu_0_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (cpu_0_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_0_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	Core3_cpu_1 cpu_1 (
		.clk                                   (clk_clk),                                                            //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                                //                   reset_n.reset_n
		.d_address                             (cpu_1_data_master_address),                                          //               data_master.address
		.d_byteenable                          (cpu_1_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (cpu_1_data_master_read),                                             //                          .read
		.d_readdata                            (cpu_1_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (cpu_1_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (cpu_1_data_master_write),                                            //                          .write
		.d_writedata                           (cpu_1_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_1_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (cpu_1_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (cpu_1_instruction_master_read),                                      //                          .read
		.i_readdata                            (cpu_1_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (cpu_1_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (cpu_1_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_1_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	Core3_onchip_memory_0 onchip_memory_0 (
		.clk        (clk_clk),                                                      //   clk1.clk
		.address    (onchip_memory_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_memory_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_memory_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_memory_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_memory_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_memory_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                               // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                            //       .reset_req
	);

	Core3_onchip_memory_1 onchip_memory_1 (
		.clk        (clk_clk),                                                      //   clk1.clk
		.address    (onchip_memory_1_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_memory_1_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_memory_1_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_memory_1_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_memory_1_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_memory_1_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory_1_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),                           // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)                        //       .reset_req
	);

	Core3_timer_0_0 timer_0_0 (
		.clk        (clk_clk),                                                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        // reset.reset_n
		.address    (timer_0_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                                //   irq.irq
	);

	Core3_timer_0_0 timer_1_0 (
		.clk        (clk_clk),                                                //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    // reset.reset_n
		.address    (timer_1_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_1_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_1_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_1_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_1_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_001_receiver0_irq)                            //   irq.irq
	);

	Core3_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                                  //               irq.irq
	);

	Core3_jtag_uart_0 jtag_uart_1 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver1_irq)                                              //               irq.irq
	);

	Core3_mutex_0 mutex_0 (
		.reset_n       (~rst_controller_002_reset_out_reset),                  // reset.reset_n
		.clk           (clk_clk),                                              //   clk.clk
		.chipselect    (mutex_0_s1_translator_avalon_anti_slave_0_chipselect), //    s1.chipselect
		.data_from_cpu (mutex_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.read          (mutex_0_s1_translator_avalon_anti_slave_0_read),       //      .read
		.write         (mutex_0_s1_translator_avalon_anti_slave_0_write),      //      .write
		.data_to_cpu   (mutex_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.address       (mutex_0_s1_translator_avalon_anti_slave_0_address)     //      .address
	);

	Core3_onchip_shared onchip_shared (
		.clk        (clk_clk),                                                    //   clk1.clk
		.address    (onchip_shared_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_shared_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_shared_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_shared_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_shared_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_shared_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_shared_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),                         // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)                      //       .reset_req
	);

	Core3_red_leds red_leds (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                   //               reset.reset_n
		.address    (red_leds_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~red_leds_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (red_leds_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (red_leds_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (red_leds_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (red_leds_external_connection_export)                    // external_connection.export
	);

	Core3_green_leds green_leds (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                     //               reset.reset_n
		.address    (green_leds_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~green_leds_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (green_leds_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (green_leds_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (green_leds_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (green_leds_external_connection_export)                    // external_connection.export
	);

	Core3_switches switches (
		.clk      (clk_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                 //               reset.reset_n
		.address  (switches_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (switches_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (switches_external_connection_export)                  // external_connection.export
	);

	Core3_fifo_0_to_1 fifo_0_to_1 (
		.wrclock                          (clk_clk),                                                      //    clk_in.clk
		.wrreset_n                        (~rst_controller_reset_out_reset),                              //  reset_in.reset_n
		.rdclock                          (clk_clk),                                                      //   clk_out.clk
		.rdreset_n                        (~rst_controller_001_reset_out_reset),                          // reset_out.reset_n
		.avalonmm_write_slave_writedata   (fifo_0_to_1_in_translator_avalon_anti_slave_0_writedata),      //        in.writedata
		.avalonmm_write_slave_write       (fifo_0_to_1_in_translator_avalon_anti_slave_0_write),          //          .write
		.avalonmm_write_slave_waitrequest (fifo_0_to_1_in_translator_avalon_anti_slave_0_waitrequest),    //          .waitrequest
		.avalonmm_read_slave_readdata     (fifo_0_to_1_out_translator_avalon_anti_slave_0_readdata),      //       out.readdata
		.avalonmm_read_slave_read         (fifo_0_to_1_out_translator_avalon_anti_slave_0_read),          //          .read
		.avalonmm_read_slave_waitrequest  (fifo_0_to_1_out_translator_avalon_anti_slave_0_waitrequest),   //          .waitrequest
		.rdclk_control_slave_address      (fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_address),   //   out_csr.address
		.rdclk_control_slave_read         (fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_read),      //          .read
		.rdclk_control_slave_writedata    (fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_writedata), //          .writedata
		.rdclk_control_slave_write        (fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_write),     //          .write
		.rdclk_control_slave_readdata     (fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_readdata),  //          .readdata
		.wrclk_control_slave_address      (fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_address),    //    in_csr.address
		.wrclk_control_slave_read         (fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_read),       //          .read
		.wrclk_control_slave_writedata    (fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_writedata),  //          .writedata
		.wrclk_control_slave_write        (fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_write),      //          .write
		.wrclk_control_slave_readdata     (fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_readdata)    //          .readdata
	);

	Core3_fifo_0_to_1 fifo_0_to_2 (
		.wrclock                          (clk_clk),                                                      //    clk_in.clk
		.wrreset_n                        (~rst_controller_reset_out_reset),                              //  reset_in.reset_n
		.rdclock                          (clk_clk),                                                      //   clk_out.clk
		.rdreset_n                        (~rst_controller_003_reset_out_reset),                          // reset_out.reset_n
		.avalonmm_write_slave_writedata   (fifo_0_to_2_in_translator_avalon_anti_slave_0_writedata),      //        in.writedata
		.avalonmm_write_slave_write       (fifo_0_to_2_in_translator_avalon_anti_slave_0_write),          //          .write
		.avalonmm_write_slave_waitrequest (fifo_0_to_2_in_translator_avalon_anti_slave_0_waitrequest),    //          .waitrequest
		.avalonmm_read_slave_readdata     (fifo_0_to_2_out_translator_avalon_anti_slave_0_readdata),      //       out.readdata
		.avalonmm_read_slave_read         (fifo_0_to_2_out_translator_avalon_anti_slave_0_read),          //          .read
		.avalonmm_read_slave_waitrequest  (fifo_0_to_2_out_translator_avalon_anti_slave_0_waitrequest),   //          .waitrequest
		.rdclk_control_slave_address      (fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_address),   //   out_csr.address
		.rdclk_control_slave_read         (fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_read),      //          .read
		.rdclk_control_slave_writedata    (fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_writedata), //          .writedata
		.rdclk_control_slave_write        (fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_write),     //          .write
		.rdclk_control_slave_readdata     (fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_readdata),  //          .readdata
		.wrclk_control_slave_address      (fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_address),    //    in_csr.address
		.wrclk_control_slave_read         (fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_read),       //          .read
		.wrclk_control_slave_writedata    (fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_writedata),  //          .writedata
		.wrclk_control_slave_write        (fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_write),      //          .write
		.wrclk_control_slave_readdata     (fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_readdata)    //          .readdata
	);

	Core3_fifo_0_to_1 fifo_1_to_0 (
		.wrclock                          (clk_clk),                                                      //    clk_in.clk
		.wrreset_n                        (~rst_controller_001_reset_out_reset),                          //  reset_in.reset_n
		.rdclock                          (clk_clk),                                                      //   clk_out.clk
		.rdreset_n                        (~rst_controller_reset_out_reset),                              // reset_out.reset_n
		.avalonmm_write_slave_writedata   (fifo_1_to_0_in_translator_avalon_anti_slave_0_writedata),      //        in.writedata
		.avalonmm_write_slave_write       (fifo_1_to_0_in_translator_avalon_anti_slave_0_write),          //          .write
		.avalonmm_write_slave_waitrequest (fifo_1_to_0_in_translator_avalon_anti_slave_0_waitrequest),    //          .waitrequest
		.avalonmm_read_slave_readdata     (fifo_1_to_0_out_translator_avalon_anti_slave_0_readdata),      //       out.readdata
		.avalonmm_read_slave_read         (fifo_1_to_0_out_translator_avalon_anti_slave_0_read),          //          .read
		.avalonmm_read_slave_waitrequest  (fifo_1_to_0_out_translator_avalon_anti_slave_0_waitrequest),   //          .waitrequest
		.rdclk_control_slave_address      (fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_address),   //   out_csr.address
		.rdclk_control_slave_read         (fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_read),      //          .read
		.rdclk_control_slave_writedata    (fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_writedata), //          .writedata
		.rdclk_control_slave_write        (fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_write),     //          .write
		.rdclk_control_slave_readdata     (fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_readdata),  //          .readdata
		.wrclk_control_slave_address      (fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_address),    //    in_csr.address
		.wrclk_control_slave_read         (fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_read),       //          .read
		.wrclk_control_slave_writedata    (fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_writedata),  //          .writedata
		.wrclk_control_slave_write        (fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_write),      //          .write
		.wrclk_control_slave_readdata     (fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_readdata)    //          .readdata
	);

	Core3_fifo_0_to_1 fifo_1_to_2 (
		.wrclock                          (clk_clk),                                                      //    clk_in.clk
		.wrreset_n                        (~rst_controller_001_reset_out_reset),                          //  reset_in.reset_n
		.rdclock                          (clk_clk),                                                      //   clk_out.clk
		.rdreset_n                        (~rst_controller_003_reset_out_reset),                          // reset_out.reset_n
		.avalonmm_write_slave_writedata   (fifo_1_to_2_in_translator_avalon_anti_slave_0_writedata),      //        in.writedata
		.avalonmm_write_slave_write       (fifo_1_to_2_in_translator_avalon_anti_slave_0_write),          //          .write
		.avalonmm_write_slave_waitrequest (fifo_1_to_2_in_translator_avalon_anti_slave_0_waitrequest),    //          .waitrequest
		.avalonmm_read_slave_readdata     (fifo_1_to_2_out_translator_avalon_anti_slave_0_readdata),      //       out.readdata
		.avalonmm_read_slave_read         (fifo_1_to_2_out_translator_avalon_anti_slave_0_read),          //          .read
		.avalonmm_read_slave_waitrequest  (fifo_1_to_2_out_translator_avalon_anti_slave_0_waitrequest),   //          .waitrequest
		.rdclk_control_slave_address      (fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_address),   //   out_csr.address
		.rdclk_control_slave_read         (fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_read),      //          .read
		.rdclk_control_slave_writedata    (fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_writedata), //          .writedata
		.rdclk_control_slave_write        (fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_write),     //          .write
		.rdclk_control_slave_readdata     (fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_readdata),  //          .readdata
		.wrclk_control_slave_address      (fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_address),    //    in_csr.address
		.wrclk_control_slave_read         (fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_read),       //          .read
		.wrclk_control_slave_writedata    (fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_writedata),  //          .writedata
		.wrclk_control_slave_write        (fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_write),      //          .write
		.wrclk_control_slave_readdata     (fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_readdata)    //          .readdata
	);

	Core3_fifo_0_to_1 fifo_2_to_0 (
		.wrclock                          (clk_clk),                                                      //    clk_in.clk
		.wrreset_n                        (~rst_controller_003_reset_out_reset),                          //  reset_in.reset_n
		.rdclock                          (clk_clk),                                                      //   clk_out.clk
		.rdreset_n                        (~rst_controller_reset_out_reset),                              // reset_out.reset_n
		.avalonmm_write_slave_writedata   (fifo_2_to_0_in_translator_avalon_anti_slave_0_writedata),      //        in.writedata
		.avalonmm_write_slave_write       (fifo_2_to_0_in_translator_avalon_anti_slave_0_write),          //          .write
		.avalonmm_write_slave_waitrequest (fifo_2_to_0_in_translator_avalon_anti_slave_0_waitrequest),    //          .waitrequest
		.avalonmm_read_slave_readdata     (fifo_2_to_0_out_translator_avalon_anti_slave_0_readdata),      //       out.readdata
		.avalonmm_read_slave_read         (fifo_2_to_0_out_translator_avalon_anti_slave_0_read),          //          .read
		.avalonmm_read_slave_waitrequest  (fifo_2_to_0_out_translator_avalon_anti_slave_0_waitrequest),   //          .waitrequest
		.rdclk_control_slave_address      (fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_address),   //   out_csr.address
		.rdclk_control_slave_read         (fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_read),      //          .read
		.rdclk_control_slave_writedata    (fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_writedata), //          .writedata
		.rdclk_control_slave_write        (fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_write),     //          .write
		.rdclk_control_slave_readdata     (fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_readdata),  //          .readdata
		.wrclk_control_slave_address      (fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_address),    //    in_csr.address
		.wrclk_control_slave_read         (fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_read),       //          .read
		.wrclk_control_slave_writedata    (fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_writedata),  //          .writedata
		.wrclk_control_slave_write        (fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_write),      //          .write
		.wrclk_control_slave_readdata     (fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_readdata)    //          .readdata
	);

	Core3_fifo_0_to_1 fifo_2_to_1 (
		.wrclock                          (clk_clk),                                                      //    clk_in.clk
		.wrreset_n                        (~rst_controller_003_reset_out_reset),                          //  reset_in.reset_n
		.rdclock                          (clk_clk),                                                      //   clk_out.clk
		.rdreset_n                        (~rst_controller_001_reset_out_reset),                          // reset_out.reset_n
		.avalonmm_write_slave_writedata   (fifo_2_to_1_in_translator_avalon_anti_slave_0_writedata),      //        in.writedata
		.avalonmm_write_slave_write       (fifo_2_to_1_in_translator_avalon_anti_slave_0_write),          //          .write
		.avalonmm_write_slave_waitrequest (fifo_2_to_1_in_translator_avalon_anti_slave_0_waitrequest),    //          .waitrequest
		.avalonmm_read_slave_readdata     (fifo_2_to_1_out_translator_avalon_anti_slave_0_readdata),      //       out.readdata
		.avalonmm_read_slave_read         (fifo_2_to_1_out_translator_avalon_anti_slave_0_read),          //          .read
		.avalonmm_read_slave_waitrequest  (fifo_2_to_1_out_translator_avalon_anti_slave_0_waitrequest),   //          .waitrequest
		.rdclk_control_slave_address      (fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_address),   //   out_csr.address
		.rdclk_control_slave_read         (fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_read),      //          .read
		.rdclk_control_slave_writedata    (fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_writedata), //          .writedata
		.rdclk_control_slave_write        (fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_write),     //          .write
		.rdclk_control_slave_readdata     (fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_readdata),  //          .readdata
		.wrclk_control_slave_address      (fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_address),    //    in_csr.address
		.wrclk_control_slave_read         (fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_read),       //          .read
		.wrclk_control_slave_writedata    (fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_writedata),  //          .writedata
		.wrclk_control_slave_write        (fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_write),      //          .write
		.wrclk_control_slave_readdata     (fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_readdata)    //          .readdata
	);

	Core3_mutex_0 mutex_1 (
		.reset_n       (~rst_controller_002_reset_out_reset),                  // reset.reset_n
		.clk           (clk_clk),                                              //   clk.clk
		.chipselect    (mutex_1_s1_translator_avalon_anti_slave_0_chipselect), //    s1.chipselect
		.data_from_cpu (mutex_1_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.read          (mutex_1_s1_translator_avalon_anti_slave_0_read),       //      .read
		.write         (mutex_1_s1_translator_avalon_anti_slave_0_write),      //      .write
		.data_to_cpu   (mutex_1_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.address       (mutex_1_s1_translator_avalon_anti_slave_0_address)     //      .address
	);

	Core3_mutex_0 mutex_2 (
		.reset_n       (~rst_controller_002_reset_out_reset),                  // reset.reset_n
		.clk           (clk_clk),                                              //   clk.clk
		.chipselect    (mutex_2_s1_translator_avalon_anti_slave_0_chipselect), //    s1.chipselect
		.data_from_cpu (mutex_2_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.read          (mutex_2_s1_translator_avalon_anti_slave_0_read),       //      .read
		.write         (mutex_2_s1_translator_avalon_anti_slave_0_write),      //      .write
		.data_to_cpu   (mutex_2_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.address       (mutex_2_s1_translator_avalon_anti_slave_0_address)     //      .address
	);

	Core3_mutex_0 mutex_3 (
		.reset_n       (~rst_controller_002_reset_out_reset),                  // reset.reset_n
		.clk           (clk_clk),                                              //   clk.clk
		.chipselect    (mutex_3_s1_translator_avalon_anti_slave_0_chipselect), //    s1.chipselect
		.data_from_cpu (mutex_3_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.read          (mutex_3_s1_translator_avalon_anti_slave_0_read),       //      .read
		.write         (mutex_3_s1_translator_avalon_anti_slave_0_write),      //      .write
		.data_to_cpu   (mutex_3_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.address       (mutex_3_s1_translator_avalon_anti_slave_0_address)     //      .address
	);

	Core3_mutex_0 mutex_4 (
		.reset_n       (~rst_controller_002_reset_out_reset),                  // reset.reset_n
		.clk           (clk_clk),                                              //   clk.clk
		.chipselect    (mutex_4_s1_translator_avalon_anti_slave_0_chipselect), //    s1.chipselect
		.data_from_cpu (mutex_4_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.read          (mutex_4_s1_translator_avalon_anti_slave_0_read),       //      .read
		.write         (mutex_4_s1_translator_avalon_anti_slave_0_write),      //      .write
		.data_to_cpu   (mutex_4_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.address       (mutex_4_s1_translator_avalon_anti_slave_0_address)     //      .address
	);

	Core3_mutex_0 mutex_5 (
		.reset_n       (~rst_controller_002_reset_out_reset),                  // reset.reset_n
		.clk           (clk_clk),                                              //   clk.clk
		.chipselect    (mutex_5_s1_translator_avalon_anti_slave_0_chipselect), //    s1.chipselect
		.data_from_cpu (mutex_5_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.read          (mutex_5_s1_translator_avalon_anti_slave_0_read),       //      .read
		.write         (mutex_5_s1_translator_avalon_anti_slave_0_write),      //      .write
		.data_to_cpu   (mutex_5_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.address       (mutex_5_s1_translator_avalon_anti_slave_0_address)     //      .address
	);

	Core3_timer_0_0 timer_shared_0 (
		.clk        (clk_clk),                                                     //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                         // reset.reset_n
		.address    (timer_shared_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_shared_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_shared_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_shared_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_shared_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                                     //   irq.irq
	);

	Core3_cpu_2 cpu_2 (
		.clk                                   (clk_clk),                                                            //                       clk.clk
		.reset_n                               (~rst_controller_003_reset_out_reset),                                //                   reset_n.reset_n
		.d_address                             (cpu_2_data_master_address),                                          //               data_master.address
		.d_byteenable                          (cpu_2_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (cpu_2_data_master_read),                                             //                          .read
		.d_readdata                            (cpu_2_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (cpu_2_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (cpu_2_data_master_write),                                            //                          .write
		.d_writedata                           (cpu_2_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_2_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (cpu_2_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (cpu_2_instruction_master_read),                                      //                          .read
		.i_readdata                            (cpu_2_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (cpu_2_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (cpu_2_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_2_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	Core3_onchip_memory_2 onchip_memory_2 (
		.clk        (clk_clk),                                                      //   clk1.clk
		.address    (onchip_memory_2_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_memory_2_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_memory_2_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_memory_2_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_memory_2_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_memory_2_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory_2_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_003_reset_out_reset),                           // reset1.reset
		.reset_req  (rst_controller_003_reset_out_reset_req)                        //       .reset_req
	);

	Core3_timer_0_0 timer_2_0 (
		.clk        (clk_clk),                                                //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                    // reset.reset_n
		.address    (timer_2_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_2_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_2_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_2_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_2_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_002_receiver0_irq)                            //   irq.irq
	);

	Core3_jtag_uart_0 jtag_uart_2 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_003_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_002_receiver1_irq)                                              //               irq.irq
	);

	Core3_performance_counter_0 performance_counter_0 (
		.clk           (clk_clk),                                                                          //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                                  //         reset.reset_n
		.address       (performance_counter_0_control_slave_translator_avalon_anti_slave_0_address),       // control_slave.address
		.begintransfer (performance_counter_0_control_slave_translator_avalon_anti_slave_0_begintransfer), //              .begintransfer
		.readdata      (performance_counter_0_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.write         (performance_counter_0_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.writedata     (performance_counter_0_control_slave_translator_avalon_anti_slave_0_writedata)      //              .writedata
	);

	Core3_performance_counter_0 performance_counter_1 (
		.clk           (clk_clk),                                                                          //           clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                                              //         reset.reset_n
		.address       (performance_counter_1_control_slave_translator_avalon_anti_slave_0_address),       // control_slave.address
		.begintransfer (performance_counter_1_control_slave_translator_avalon_anti_slave_0_begintransfer), //              .begintransfer
		.readdata      (performance_counter_1_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.write         (performance_counter_1_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.writedata     (performance_counter_1_control_slave_translator_avalon_anti_slave_0_writedata)      //              .writedata
	);

	Core3_performance_counter_0 performance_counter_2 (
		.clk           (clk_clk),                                                                          //           clk.clk
		.reset_n       (~rst_controller_003_reset_out_reset),                                              //         reset.reset_n
		.address       (performance_counter_2_control_slave_translator_avalon_anti_slave_0_address),       // control_slave.address
		.begintransfer (performance_counter_2_control_slave_translator_avalon_anti_slave_0_begintransfer), //              .begintransfer
		.readdata      (performance_counter_2_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.write         (performance_counter_2_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.writedata     (performance_counter_2_control_slave_translator_avalon_anti_slave_0_writedata)      //              .writedata
	);

	Core3_timer_0_0 timer_0_1 (
		.clk        (clk_clk),                                                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        // reset.reset_n
		.address    (timer_0_1_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_1_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_1_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_1_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_1_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                                //   irq.irq
	);

	Core3_timer_0_0 timer_1_1 (
		.clk        (clk_clk),                                                //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    // reset.reset_n
		.address    (timer_1_1_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_1_1_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_1_1_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_1_1_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_1_1_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_001_receiver3_irq)                            //   irq.irq
	);

	Core3_timer_0_0 timer_2_1 (
		.clk        (clk_clk),                                                //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                    // reset.reset_n
		.address    (timer_2_1_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_2_1_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_2_1_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_2_1_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_2_1_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_002_receiver3_irq)                            //   irq.irq
	);

	Core3_timer_0_0 timer_shared_1 (
		.clk        (clk_clk),                                                     //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                         // reset.reset_n
		.address    (timer_shared_1_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_shared_1_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_shared_1_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_shared_1_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_shared_1_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                                     //   irq.irq
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (18),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (18),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_0_instruction_master_translator (
		.clk                      (clk_clk),                                                                     //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address              (cpu_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (cpu_0_instruction_master_read),                                               //                          .read
		.av_readdata              (cpu_0_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_byteenable            (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_readdatavalid         (),                                                                            //               (terminated)
		.av_write                 (1'b0),                                                                        //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.av_debugaccess           (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (18),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (18),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) cpu_0_data_master_translator (
		.clk                      (clk_clk),                                                              //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address              (cpu_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (cpu_0_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (cpu_0_data_master_read),                                               //                          .read
		.av_readdata              (cpu_0_data_master_readdata),                                           //                          .readdata
		.av_write                 (cpu_0_data_master_write),                                              //                          .write
		.av_writedata             (cpu_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (cpu_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                 //               (terminated)
		.av_begintransfer         (1'b0),                                                                 //               (terminated)
		.av_chipselect            (1'b0),                                                                 //               (terminated)
		.av_readdatavalid         (),                                                                     //               (terminated)
		.av_lock                  (1'b0),                                                                 //               (terminated)
		.uav_clken                (),                                                                     //               (terminated)
		.av_clken                 (1'b1),                                                                 //               (terminated)
		.uav_response             (2'b00),                                                                //               (terminated)
		.av_response              (),                                                                     //               (terminated)
		.uav_writeresponserequest (),                                                                     //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                 //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                 //               (terminated)
		.av_writeresponsevalid    ()                                                                      //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (18),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (18),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) cpu_1_data_master_translator (
		.clk                      (clk_clk),                                                              //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                   //                     reset.reset
		.uav_address              (cpu_1_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_1_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_1_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_1_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_1_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_1_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_1_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_1_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_1_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_1_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_1_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_1_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_1_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (cpu_1_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (cpu_1_data_master_read),                                               //                          .read
		.av_readdata              (cpu_1_data_master_readdata),                                           //                          .readdata
		.av_write                 (cpu_1_data_master_write),                                              //                          .write
		.av_writedata             (cpu_1_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (cpu_1_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                 //               (terminated)
		.av_begintransfer         (1'b0),                                                                 //               (terminated)
		.av_chipselect            (1'b0),                                                                 //               (terminated)
		.av_readdatavalid         (),                                                                     //               (terminated)
		.av_lock                  (1'b0),                                                                 //               (terminated)
		.uav_clken                (),                                                                     //               (terminated)
		.av_clken                 (1'b1),                                                                 //               (terminated)
		.uav_response             (2'b00),                                                                //               (terminated)
		.av_response              (),                                                                     //               (terminated)
		.uav_writeresponserequest (),                                                                     //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                 //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                 //               (terminated)
		.av_writeresponsevalid    ()                                                                      //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (18),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (18),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) cpu_2_data_master_translator (
		.clk                      (clk_clk),                                                              //                       clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                   //                     reset.reset
		.uav_address              (cpu_2_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_2_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_2_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_2_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_2_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_2_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_2_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_2_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_2_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_2_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_2_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_2_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_2_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (cpu_2_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (cpu_2_data_master_read),                                               //                          .read
		.av_readdata              (cpu_2_data_master_readdata),                                           //                          .readdata
		.av_write                 (cpu_2_data_master_write),                                              //                          .write
		.av_writedata             (cpu_2_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (cpu_2_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                 //               (terminated)
		.av_begintransfer         (1'b0),                                                                 //               (terminated)
		.av_chipselect            (1'b0),                                                                 //               (terminated)
		.av_readdatavalid         (),                                                                     //               (terminated)
		.av_lock                  (1'b0),                                                                 //               (terminated)
		.uav_clken                (),                                                                     //               (terminated)
		.av_clken                 (1'b1),                                                                 //               (terminated)
		.uav_response             (2'b00),                                                                //               (terminated)
		.av_response              (),                                                                     //               (terminated)
		.uav_writeresponserequest (),                                                                     //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                 //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                 //               (terminated)
		.av_writeresponsevalid    ()                                                                      //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (18),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (18),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_1_instruction_master_translator (
		.clk                      (clk_clk),                                                                     //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                          //                     reset.reset
		.uav_address              (cpu_1_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_1_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_1_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_1_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_1_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_1_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_1_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_1_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_1_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_1_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_1_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_1_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_1_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (cpu_1_instruction_master_read),                                               //                          .read
		.av_readdata              (cpu_1_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_byteenable            (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_readdatavalid         (),                                                                            //               (terminated)
		.av_write                 (1'b0),                                                                        //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.av_debugaccess           (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (18),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (18),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_2_instruction_master_translator (
		.clk                      (clk_clk),                                                                     //                       clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                          //                     reset.reset
		.uav_address              (cpu_2_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_2_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_2_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_2_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_2_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_2_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_2_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_2_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_2_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_2_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_2_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_2_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_2_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (cpu_2_instruction_master_read),                                               //                          .read
		.av_readdata              (cpu_2_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_byteenable            (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_readdatavalid         (),                                                                            //               (terminated)
		.av_write                 (1'b0),                                                                        //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.av_debugaccess           (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_0_jtag_debug_module_translator (
		.clk                      (clk_clk),                                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_chipselect            (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory_0_s1_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address              (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                              //              (terminated)
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (14),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_shared_s1_translator (
		.clk                      (clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                          //                    reset.reset
		.uav_address              (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_shared_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_shared_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_shared_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_shared_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_shared_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_shared_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_shared_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_0_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address              (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_0_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_0_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_0_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_0_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_0_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mutex_0_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                    //                    reset.reset
		.uav_address              (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (mutex_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (mutex_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (mutex_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (mutex_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (mutex_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (mutex_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mutex_1_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                    //                    reset.reset
		.uav_address              (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (mutex_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (mutex_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (mutex_1_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (mutex_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (mutex_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (mutex_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mutex_2_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                    //                    reset.reset
		.uav_address              (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (mutex_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (mutex_2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (mutex_2_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (mutex_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (mutex_2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (mutex_2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mutex_3_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                    //                    reset.reset
		.uav_address              (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (mutex_3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (mutex_3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (mutex_3_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (mutex_3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (mutex_3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (mutex_3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mutex_4_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                    //                    reset.reset
		.uav_address              (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (mutex_4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (mutex_4_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (mutex_4_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (mutex_4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (mutex_4_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (mutex_4_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mutex_5_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                    //                    reset.reset
		.uav_address              (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (mutex_5_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (mutex_5_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (mutex_5_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (mutex_5_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (mutex_5_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (mutex_5_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_to_1_in_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                    reset.reset
		.uav_address              (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (fifo_0_to_1_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata             (fifo_0_to_1_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (fifo_0_to_1_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address               (),                                                                          //              (terminated)
		.av_read                  (),                                                                          //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                      //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_chipselect            (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_to_1_in_csr_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address              (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_0_to_1_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_chipselect            (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_to_2_in_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                    reset.reset
		.uav_address              (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (fifo_0_to_2_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata             (fifo_0_to_2_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (fifo_0_to_2_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address               (),                                                                          //              (terminated)
		.av_read                  (),                                                                          //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                      //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_chipselect            (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_to_2_in_csr_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address              (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_0_to_2_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_chipselect            (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_1_to_0_out_csr_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_1_to_0_out_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_1_to_0_out_translator (
		.clk                      (clk_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                             //                    reset.reset
		.uav_address              (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read                  (fifo_1_to_0_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata              (fifo_1_to_0_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest           (fifo_1_to_0_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address               (),                                                                           //              (terminated)
		.av_write                 (),                                                                           //              (terminated)
		.av_writedata             (),                                                                           //              (terminated)
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_chipselect            (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_2_to_0_out_translator (
		.clk                      (clk_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                             //                    reset.reset
		.uav_address              (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read                  (fifo_2_to_0_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata              (fifo_2_to_0_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest           (fifo_2_to_0_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address               (),                                                                           //              (terminated)
		.av_write                 (),                                                                           //              (terminated)
		.av_writedata             (),                                                                           //              (terminated)
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_chipselect            (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_2_to_0_out_csr_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_2_to_0_out_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) red_leds_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                     //                    reset.reset
		.uav_address              (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (red_leds_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (red_leds_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (red_leds_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (red_leds_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (red_leds_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) green_leds_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                       //                    reset.reset
		.uav_address              (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (green_leds_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (green_leds_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (green_leds_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (green_leds_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (green_leds_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switches_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                     //                    reset.reset
		.uav_address              (switches_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switches_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switches_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (switches_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                       //              (terminated)
		.av_read                  (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_shared_0_s1_translator (
		.clk                      (clk_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                           //                    reset.reset
		.uav_address              (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_shared_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_shared_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_shared_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_shared_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_shared_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (5),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) performance_counter_0_control_slave_translator (
		.clk                      (clk_clk),                                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                 //                    reset.reset
		.uav_address              (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (performance_counter_0_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (performance_counter_0_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (performance_counter_0_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (performance_counter_0_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (performance_counter_0_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_read                  (),                                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                                               //              (terminated)
		.av_burstcount            (),                                                                                               //              (terminated)
		.av_byteenable            (),                                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                                               //              (terminated)
		.av_lock                  (),                                                                                               //              (terminated)
		.av_chipselect            (),                                                                                               //              (terminated)
		.av_clken                 (),                                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                                           //              (terminated)
		.av_debugaccess           (),                                                                                               //              (terminated)
		.av_outputenable          (),                                                                                               //              (terminated)
		.uav_response             (),                                                                                               //              (terminated)
		.av_response              (2'b00),                                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_1_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address              (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_0_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_0_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_0_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_0_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_0_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_shared_1_s1_translator (
		.clk                      (clk_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                           //                    reset.reset
		.uav_address              (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_shared_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_shared_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_shared_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_shared_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_shared_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_1_jtag_debug_module_translator (
		.clk                      (clk_clk),                                                                            //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (cpu_1_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_chipselect            (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory_1_s1_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                            //                    reset.reset
		.uav_address              (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory_1_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory_1_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                              //              (terminated)
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_1_0_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_1_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_1_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_1_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_1_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_1_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_1_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                       //                    reset.reset
		.uav_address              (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_1_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_to_1_out_translator (
		.clk                      (clk_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                         //                    reset.reset
		.uav_address              (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read                  (fifo_0_to_1_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata              (fifo_0_to_1_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest           (fifo_0_to_1_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address               (),                                                                           //              (terminated)
		.av_write                 (),                                                                           //              (terminated)
		.av_writedata             (),                                                                           //              (terminated)
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_chipselect            (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_to_1_out_csr_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                             //                    reset.reset
		.uav_address              (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_0_to_1_out_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_1_to_0_in_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (fifo_1_to_0_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata             (fifo_1_to_0_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (fifo_1_to_0_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address               (),                                                                          //              (terminated)
		.av_read                  (),                                                                          //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                      //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_chipselect            (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_1_to_0_in_csr_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                            //                    reset.reset
		.uav_address              (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_1_to_0_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_chipselect            (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_1_to_2_in_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (fifo_1_to_2_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata             (fifo_1_to_2_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (fifo_1_to_2_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address               (),                                                                          //              (terminated)
		.av_read                  (),                                                                          //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                      //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_chipselect            (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_1_to_2_in_csr_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                            //                    reset.reset
		.uav_address              (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_1_to_2_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_chipselect            (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_2_to_1_out_translator (
		.clk                      (clk_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                         //                    reset.reset
		.uav_address              (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read                  (fifo_2_to_1_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata              (fifo_2_to_1_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest           (fifo_2_to_1_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address               (),                                                                           //              (terminated)
		.av_write                 (),                                                                           //              (terminated)
		.av_writedata             (),                                                                           //              (terminated)
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_chipselect            (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_2_to_1_out_csr_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                             //                    reset.reset
		.uav_address              (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_2_to_1_out_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (5),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) performance_counter_1_control_slave_translator (
		.clk                      (clk_clk),                                                                                        //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                             //                    reset.reset
		.uav_address              (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (performance_counter_1_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (performance_counter_1_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (performance_counter_1_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (performance_counter_1_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (performance_counter_1_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_read                  (),                                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                                               //              (terminated)
		.av_burstcount            (),                                                                                               //              (terminated)
		.av_byteenable            (),                                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                                               //              (terminated)
		.av_lock                  (),                                                                                               //              (terminated)
		.av_chipselect            (),                                                                                               //              (terminated)
		.av_clken                 (),                                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                                           //              (terminated)
		.av_debugaccess           (),                                                                                               //              (terminated)
		.av_outputenable          (),                                                                                               //              (terminated)
		.uav_response             (),                                                                                               //              (terminated)
		.av_response              (2'b00),                                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_1_1_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_1_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_1_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_1_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_1_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_1_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_2_jtag_debug_module_translator (
		.clk                      (clk_clk),                                                                            //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (cpu_2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_chipselect            (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory_2_s1_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                            //                    reset.reset
		.uav_address              (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory_2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory_2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory_2_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory_2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory_2_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                              //              (terminated)
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_2_0_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                      //                    reset.reset
		.uav_address              (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_2_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_2_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_2_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_2_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_2_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_2_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                  //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                                       //                    reset.reset
		.uav_address              (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_2_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_to_2_out_translator (
		.clk                      (clk_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                         //                    reset.reset
		.uav_address              (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read                  (fifo_0_to_2_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata              (fifo_0_to_2_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest           (fifo_0_to_2_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address               (),                                                                           //              (terminated)
		.av_write                 (),                                                                           //              (terminated)
		.av_writedata             (),                                                                           //              (terminated)
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_chipselect            (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_to_2_out_csr_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                             //                    reset.reset
		.uav_address              (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_0_to_2_out_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_1_to_2_out_translator (
		.clk                      (clk_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                         //                    reset.reset
		.uav_address              (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read                  (fifo_1_to_2_out_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata              (fifo_1_to_2_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest           (fifo_1_to_2_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address               (),                                                                           //              (terminated)
		.av_write                 (),                                                                           //              (terminated)
		.av_writedata             (),                                                                           //              (terminated)
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_chipselect            (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_1_to_2_out_csr_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                             //                    reset.reset
		.uav_address              (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_1_to_2_out_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_2_to_0_in_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                        //                    reset.reset
		.uav_address              (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (fifo_2_to_0_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata             (fifo_2_to_0_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (fifo_2_to_0_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address               (),                                                                          //              (terminated)
		.av_read                  (),                                                                          //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                      //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_chipselect            (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_2_to_0_in_csr_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                            //                    reset.reset
		.uav_address              (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_2_to_0_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_chipselect            (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_2_to_1_in_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                        //                    reset.reset
		.uav_address              (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (fifo_2_to_1_in_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata             (fifo_2_to_1_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (fifo_2_to_1_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address               (),                                                                          //              (terminated)
		.av_read                  (),                                                                          //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                      //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_chipselect            (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_2_to_1_in_csr_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                            //                    reset.reset
		.uav_address              (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_2_to_1_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_chipselect            (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (5),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) performance_counter_2_control_slave_translator (
		.clk                      (clk_clk),                                                                                        //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                                             //                    reset.reset
		.uav_address              (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (performance_counter_2_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (performance_counter_2_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (performance_counter_2_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (performance_counter_2_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (performance_counter_2_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_read                  (),                                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                                               //              (terminated)
		.av_burstcount            (),                                                                                               //              (terminated)
		.av_byteenable            (),                                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                                               //              (terminated)
		.av_lock                  (),                                                                                               //              (terminated)
		.av_chipselect            (),                                                                                               //              (terminated)
		.av_clken                 (),                                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                                           //              (terminated)
		.av_debugaccess           (),                                                                                               //              (terminated)
		.av_outputenable          (),                                                                                               //              (terminated)
		.uav_response             (),                                                                                               //              (terminated)
		.av_response              (2'b00),                                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_2_1_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                      //                    reset.reset
		.uav_address              (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_2_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_2_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_2_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_2_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_2_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (73),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.PKT_BURST_TYPE_H          (70),
		.PKT_BURST_TYPE_L          (69),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_TRANS_EXCLUSIVE       (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_THREAD_ID_H           (87),
		.PKT_THREAD_ID_L           (87),
		.PKT_CACHE_H               (94),
		.PKT_CACHE_L               (91),
		.PKT_DATA_SIDEBAND_H       (72),
		.PKT_DATA_SIDEBAND_L       (72),
		.PKT_QOS_H                 (74),
		.PKT_QOS_L                 (74),
		.PKT_ADDR_SIDEBAND_H       (71),
		.PKT_ADDR_SIDEBAND_L       (71),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.ST_DATA_W                 (97),
		.ST_CHANNEL_W              (54),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                              //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address              (cpu_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                               //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                             //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                       //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                         //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                               //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (73),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.PKT_BURST_TYPE_H          (70),
		.PKT_BURST_TYPE_L          (69),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_TRANS_EXCLUSIVE       (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_THREAD_ID_H           (87),
		.PKT_THREAD_ID_L           (87),
		.PKT_CACHE_H               (94),
		.PKT_CACHE_L               (91),
		.PKT_DATA_SIDEBAND_H       (72),
		.PKT_DATA_SIDEBAND_L       (72),
		.PKT_QOS_H                 (74),
		.PKT_QOS_L                 (74),
		.PKT_ADDR_SIDEBAND_H       (71),
		.PKT_ADDR_SIDEBAND_L       (71),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.ST_DATA_W                 (97),
		.ST_CHANNEL_W              (54),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_0_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                       //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address              (cpu_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                    //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                     //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                  //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                              //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                    //          .ready
		.av_response             (),                                                                              // (terminated)
		.av_writeresponserequest (1'b0),                                                                          // (terminated)
		.av_writeresponsevalid   ()                                                                               // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (73),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.PKT_BURST_TYPE_H          (70),
		.PKT_BURST_TYPE_L          (69),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_TRANS_EXCLUSIVE       (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_THREAD_ID_H           (87),
		.PKT_THREAD_ID_L           (87),
		.PKT_CACHE_H               (94),
		.PKT_CACHE_L               (91),
		.PKT_DATA_SIDEBAND_H       (72),
		.PKT_DATA_SIDEBAND_L       (72),
		.PKT_QOS_H                 (74),
		.PKT_QOS_L                 (74),
		.PKT_ADDR_SIDEBAND_H       (71),
		.PKT_ADDR_SIDEBAND_L       (71),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.ST_DATA_W                 (97),
		.ST_CHANNEL_W              (54),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_1_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                       //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.av_address              (cpu_1_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_1_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_1_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_1_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_1_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_1_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_1_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_1_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_1_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_1_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_1_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_002_src_valid),                                                    //        rp.valid
		.rp_data                 (rsp_xbar_mux_002_src_data),                                                     //          .data
		.rp_channel              (rsp_xbar_mux_002_src_channel),                                                  //          .channel
		.rp_startofpacket        (rsp_xbar_mux_002_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_002_src_endofpacket),                                              //          .endofpacket
		.rp_ready                (rsp_xbar_mux_002_src_ready),                                                    //          .ready
		.av_response             (),                                                                              // (terminated)
		.av_writeresponserequest (1'b0),                                                                          // (terminated)
		.av_writeresponsevalid   ()                                                                               // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (73),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.PKT_BURST_TYPE_H          (70),
		.PKT_BURST_TYPE_L          (69),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_TRANS_EXCLUSIVE       (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_THREAD_ID_H           (87),
		.PKT_THREAD_ID_L           (87),
		.PKT_CACHE_H               (94),
		.PKT_CACHE_L               (91),
		.PKT_DATA_SIDEBAND_H       (72),
		.PKT_DATA_SIDEBAND_L       (72),
		.PKT_QOS_H                 (74),
		.PKT_QOS_L                 (74),
		.PKT_ADDR_SIDEBAND_H       (71),
		.PKT_ADDR_SIDEBAND_L       (71),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.ST_DATA_W                 (97),
		.ST_CHANNEL_W              (54),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_1_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                              //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.av_address              (cpu_1_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_1_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_1_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_1_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_1_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_1_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_1_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_1_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_1_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_1_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_1_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_003_src_valid),                                                           //        rp.valid
		.rp_data                 (rsp_xbar_mux_003_src_data),                                                            //          .data
		.rp_channel              (rsp_xbar_mux_003_src_channel),                                                         //          .channel
		.rp_startofpacket        (rsp_xbar_mux_003_src_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_003_src_endofpacket),                                                     //          .endofpacket
		.rp_ready                (rsp_xbar_mux_003_src_ready),                                                           //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (73),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.PKT_BURST_TYPE_H          (70),
		.PKT_BURST_TYPE_L          (69),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_TRANS_EXCLUSIVE       (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_THREAD_ID_H           (87),
		.PKT_THREAD_ID_L           (87),
		.PKT_CACHE_H               (94),
		.PKT_CACHE_L               (91),
		.PKT_DATA_SIDEBAND_H       (72),
		.PKT_DATA_SIDEBAND_L       (72),
		.PKT_QOS_H                 (74),
		.PKT_QOS_L                 (74),
		.PKT_ADDR_SIDEBAND_H       (71),
		.PKT_ADDR_SIDEBAND_L       (71),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.ST_DATA_W                 (97),
		.ST_CHANNEL_W              (54),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (4),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_2_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                       //       clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                            // clk_reset.reset
		.av_address              (cpu_2_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_2_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_2_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_2_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_2_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_2_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_2_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_2_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_2_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_2_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_2_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_004_src_valid),                                                    //        rp.valid
		.rp_data                 (rsp_xbar_mux_004_src_data),                                                     //          .data
		.rp_channel              (rsp_xbar_mux_004_src_channel),                                                  //          .channel
		.rp_startofpacket        (rsp_xbar_mux_004_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_004_src_endofpacket),                                              //          .endofpacket
		.rp_ready                (rsp_xbar_mux_004_src_ready),                                                    //          .ready
		.av_response             (),                                                                              // (terminated)
		.av_writeresponserequest (1'b0),                                                                          // (terminated)
		.av_writeresponsevalid   ()                                                                               // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (73),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.PKT_BURST_TYPE_H          (70),
		.PKT_BURST_TYPE_L          (69),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_TRANS_EXCLUSIVE       (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_THREAD_ID_H           (87),
		.PKT_THREAD_ID_L           (87),
		.PKT_CACHE_H               (94),
		.PKT_CACHE_L               (91),
		.PKT_DATA_SIDEBAND_H       (72),
		.PKT_DATA_SIDEBAND_L       (72),
		.PKT_QOS_H                 (74),
		.PKT_QOS_L                 (74),
		.PKT_ADDR_SIDEBAND_H       (71),
		.PKT_ADDR_SIDEBAND_L       (71),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.ST_DATA_W                 (97),
		.ST_CHANNEL_W              (54),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (5),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_2_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                              //       clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.av_address              (cpu_2_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_2_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_2_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_2_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_2_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_2_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_2_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_2_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_2_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_2_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_2_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_005_src_valid),                                                           //        rp.valid
		.rp_data                 (rsp_xbar_mux_005_src_data),                                                            //          .data
		.rp_channel              (rsp_xbar_mux_005_src_channel),                                                         //          .channel
		.rp_startofpacket        (rsp_xbar_mux_005_src_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_005_src_endofpacket),                                                     //          .endofpacket
		.rp_ready                (rsp_xbar_mux_005_src_ready),                                                           //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                     //                .channel
		.rf_sink_ready           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                            //                .channel
		.rf_sink_ready           (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_shared_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_shared_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                          //                .channel
		.rf_sink_ready           (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_0_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                   //                .channel
		.rf_sink_ready           (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) mutex_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mutex_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_005_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_005_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_005_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_005_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_005_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_005_src_channel),                                                    //                .channel
		.rf_sink_ready           (mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mutex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mutex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (mutex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (mutex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mutex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mutex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.in_data           (mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mutex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mutex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) mutex_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mutex_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_006_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_006_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_006_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_006_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_006_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_006_src_channel),                                                    //                .channel
		.rf_sink_ready           (mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mutex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mutex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (mutex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (mutex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mutex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mutex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.in_data           (mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mutex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mutex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) mutex_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mutex_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_007_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_007_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_007_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_007_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_007_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_007_src_channel),                                                    //                .channel
		.rf_sink_ready           (mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mutex_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mutex_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (mutex_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (mutex_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mutex_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mutex_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.in_data           (mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mutex_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mutex_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) mutex_3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mutex_3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_008_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_008_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_008_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_008_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_008_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_008_src_channel),                                                    //                .channel
		.rf_sink_ready           (mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mutex_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mutex_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (mutex_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (mutex_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mutex_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mutex_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.in_data           (mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mutex_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mutex_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) mutex_4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mutex_4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_009_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_009_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_009_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_009_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_009_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_009_src_channel),                                                    //                .channel
		.rf_sink_ready           (mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mutex_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mutex_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (mutex_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (mutex_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mutex_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mutex_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.in_data           (mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mutex_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mutex_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) mutex_5_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mutex_5_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_010_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_010_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_010_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_010_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_010_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_010_src_channel),                                                    //                .channel
		.rf_sink_ready           (mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mutex_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mutex_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (mutex_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (mutex_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mutex_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mutex_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.in_data           (mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mutex_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mutex_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_0_to_1_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                    //                .channel
		.rf_sink_ready           (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                        //                .channel
		.rf_sink_ready           (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_0_to_2_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src13_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src13_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src13_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src13_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src13_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src13_channel),                                                    //                .channel
		.rf_sink_ready           (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src14_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src14_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_001_src14_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src14_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src14_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src14_channel),                                                        //                .channel
		.rf_sink_ready           (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src15_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src15_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_001_src15_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src15_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src15_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src15_channel),                                                         //                .channel
		.rf_sink_ready           (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_1_to_0_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src16_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src16_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src16_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src16_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src16_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src16_channel),                                                     //                .channel
		.rf_sink_ready           (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_2_to_0_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src17_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src17_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src17_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src17_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src17_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src17_channel),                                                     //                .channel
		.rf_sink_ready           (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src18_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src18_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_001_src18_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src18_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src18_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src18_channel),                                                         //                .channel
		.rf_sink_ready           (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) red_leds_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (red_leds_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_019_src_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_019_src_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_019_src_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_019_src_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_019_src_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_019_src_channel),                                                     //                .channel
		.rf_sink_ready           (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                               // clk_reset.reset
		.in_data           (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) green_leds_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_020_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_020_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_020_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_020_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_020_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_020_src_channel),                                                       //                .channel
		.rf_sink_ready           (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switches_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (switches_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switches_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switches_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switches_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switches_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_021_src_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_021_src_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_021_src_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_021_src_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_021_src_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_021_src_channel),                                                     //                .channel
		.rf_sink_ready           (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                               // clk_reset.reset
		.in_data           (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_shared_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_022_src_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_mux_022_src_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_mux_022_src_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_mux_022_src_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_022_src_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_mux_022_src_channel),                                                           //                .channel
		.rf_sink_ready           (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                           //       clk_reset.reset
		.m0_address              (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src23_ready),                                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src23_valid),                                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_001_src23_data),                                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src23_startofpacket),                                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src23_endofpacket),                                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src23_channel),                                                                         //                .channel
		.rf_sink_ready           (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                           // clk_reset.reset
		.in_data           (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                                     // (terminated)
		.csr_readdata      (),                                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                     // (terminated)
		.almost_full_data  (),                                                                                                         // (terminated)
		.almost_empty_data (),                                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                                     // (terminated)
		.out_empty         (),                                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                                     // (terminated)
		.out_error         (),                                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                                     // (terminated)
		.out_channel       ()                                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_0_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src24_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src24_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src24_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src24_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src24_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src24_channel),                                                  //                .channel
		.rf_sink_ready           (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_shared_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_025_src_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_mux_025_src_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_mux_025_src_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_mux_025_src_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_025_src_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_mux_025_src_channel),                                                           //                .channel
		.rf_sink_ready           (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_026_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_026_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_026_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_026_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_026_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_026_src_channel),                                                                 //                .channel
		.rf_sink_ready           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_027_src_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_027_src_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_027_src_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_027_src_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_027_src_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_027_src_channel),                                                            //                .channel
		.rf_sink_ready           (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_1_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_1_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src14_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src14_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_002_src14_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src14_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src14_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src14_channel),                                                  //                .channel
		.rf_sink_ready           (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src15_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src15_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_002_src15_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src15_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src15_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src15_channel),                                                                   //                .channel
		.rf_sink_ready           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_0_to_1_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src16_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src16_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_002_src16_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src16_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src16_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src16_channel),                                                     //                .channel
		.rf_sink_ready           (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src17_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src17_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_002_src17_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src17_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src17_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src17_channel),                                                         //                .channel
		.rf_sink_ready           (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_1_to_0_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src18_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src18_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_002_src18_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src18_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src18_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src18_channel),                                                    //                .channel
		.rf_sink_ready           (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src19_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src19_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_002_src19_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src19_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src19_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src19_channel),                                                        //                .channel
		.rf_sink_ready           (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_1_to_2_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src20_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src20_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_002_src20_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src20_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src20_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src20_channel),                                                    //                .channel
		.rf_sink_ready           (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src21_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src21_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_002_src21_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src21_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src21_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src21_channel),                                                        //                .channel
		.rf_sink_ready           (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_2_to_1_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src22_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src22_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_002_src22_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src22_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src22_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src22_channel),                                                     //                .channel
		.rf_sink_ready           (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src23_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src23_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_002_src23_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src23_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src23_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src23_channel),                                                         //                .channel
		.rf_sink_ready           (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                       //       clk_reset.reset
		.m0_address              (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src24_ready),                                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src24_valid),                                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_002_src24_data),                                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src24_startofpacket),                                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src24_endofpacket),                                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src24_channel),                                                                         //                .channel
		.rf_sink_ready           (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                       // clk_reset.reset
		.in_data           (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                                     // (terminated)
		.csr_readdata      (),                                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                     // (terminated)
		.almost_full_data  (),                                                                                                         // (terminated)
		.almost_empty_data (),                                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                                     // (terminated)
		.out_empty         (),                                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                                     // (terminated)
		.out_error         (),                                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                                     // (terminated)
		.out_channel       ()                                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_1_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_1_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src25_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src25_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_002_src25_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src25_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src25_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src25_channel),                                                  //                .channel
		.rf_sink_ready           (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_040_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_040_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_040_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_040_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_040_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_040_src_channel),                                                                 //                .channel
		.rf_sink_ready           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_041_src_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_041_src_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_041_src_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_041_src_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_041_src_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_041_src_channel),                                                            //                .channel
		.rf_sink_ready           (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_2_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src14_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src14_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_004_src14_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src14_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src14_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src14_channel),                                                  //                .channel
		.rf_sink_ready           (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                // clk_reset.reset
		.in_data           (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src15_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src15_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_004_src15_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src15_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src15_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src15_channel),                                                                   //                .channel
		.rf_sink_ready           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_0_to_2_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src16_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src16_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_004_src16_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src16_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src16_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src16_channel),                                                     //                .channel
		.rf_sink_ready           (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src17_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src17_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_004_src17_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src17_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src17_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src17_channel),                                                         //                .channel
		.rf_sink_ready           (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_1_to_2_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src18_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src18_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_004_src18_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src18_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src18_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src18_channel),                                                     //                .channel
		.rf_sink_ready           (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src19_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src19_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_004_src19_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src19_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src19_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src19_channel),                                                         //                .channel
		.rf_sink_ready           (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_2_to_0_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src20_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src20_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_004_src20_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src20_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src20_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src20_channel),                                                    //                .channel
		.rf_sink_ready           (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src21_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src21_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_004_src21_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src21_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src21_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src21_channel),                                                        //                .channel
		.rf_sink_ready           (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_2_to_1_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src22_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src22_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_004_src22_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src22_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src22_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src22_channel),                                                    //                .channel
		.rf_sink_ready           (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src23_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src23_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_004_src23_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src23_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src23_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src23_channel),                                                        //                .channel
		.rf_sink_ready           (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                  //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                                       //       clk_reset.reset
		.m0_address              (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src24_ready),                                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src24_valid),                                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_004_src24_data),                                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src24_startofpacket),                                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src24_endofpacket),                                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src24_channel),                                                                         //                .channel
		.rf_sink_ready           (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                  //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                                       // clk_reset.reset
		.in_data           (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                                     // (terminated)
		.csr_readdata      (),                                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                     // (terminated)
		.almost_full_data  (),                                                                                                         // (terminated)
		.almost_empty_data (),                                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                                     // (terminated)
		.out_empty         (),                                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                                     // (terminated)
		.out_error         (),                                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                                     // (terminated)
		.out_channel       ()                                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (90),
		.PKT_PROTECTION_L          (88),
		.PKT_RESPONSE_STATUS_H     (96),
		.PKT_RESPONSE_STATUS_L     (95),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (54),
		.ST_DATA_W                 (97),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_2_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_2_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src25_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src25_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_004_src25_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src25_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src25_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src25_channel),                                                  //                .channel
		.rf_sink_ready           (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (98),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                // clk_reset.reset
		.in_data           (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	Core3_addr_router addr_router (
		.sink_ready         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_src_valid),                                                                //          .valid
		.src_data           (addr_router_src_data),                                                                 //          .data
		.src_channel        (addr_router_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                           //          .endofpacket
	);

	Core3_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                     //          .valid
		.src_data           (addr_router_001_src_data),                                                      //          .data
		.src_channel        (addr_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                //          .endofpacket
	);

	Core3_addr_router_002 addr_router_002 (
		.sink_ready         (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_1_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                     //          .valid
		.src_data           (addr_router_002_src_data),                                                      //          .data
		.src_channel        (addr_router_002_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                //          .endofpacket
	);

	Core3_addr_router_003 addr_router_003 (
		.sink_ready         (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_1_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                            //          .valid
		.src_data           (addr_router_003_src_data),                                                             //          .data
		.src_channel        (addr_router_003_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                       //          .endofpacket
	);

	Core3_addr_router_004 addr_router_004 (
		.sink_ready         (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                     //          .valid
		.src_data           (addr_router_004_src_data),                                                      //          .data
		.src_channel        (addr_router_004_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                //          .endofpacket
	);

	Core3_addr_router_005 addr_router_005 (
		.sink_ready         (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                            //          .valid
		.src_data           (addr_router_005_src_data),                                                             //          .data
		.src_channel        (addr_router_005_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                       //          .endofpacket
	);

	Core3_id_router id_router (
		.sink_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                //       src.ready
		.src_valid          (id_router_src_valid),                                                                //          .valid
		.src_data           (id_router_src_data),                                                                 //          .data
		.src_channel        (id_router_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                           //          .endofpacket
	);

	Core3_id_router id_router_001 (
		.sink_ready         (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                       //       src.ready
		.src_valid          (id_router_001_src_valid),                                                       //          .valid
		.src_data           (id_router_001_src_data),                                                        //          .data
		.src_channel        (id_router_001_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                  //          .endofpacket
	);

	Core3_id_router_002 id_router_002 (
		.sink_ready         (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_shared_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                     //       src.ready
		.src_valid          (id_router_002_src_valid),                                                     //          .valid
		.src_data           (id_router_002_src_data),                                                      //          .data
		.src_channel        (id_router_002_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                //          .endofpacket
	);

	Core3_id_router_003 id_router_003 (
		.sink_ready         (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                 //       src.ready
		.src_valid          (id_router_003_src_valid),                                                 //          .valid
		.src_data           (id_router_003_src_data),                                                  //          .data
		.src_channel        (id_router_003_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                            //          .endofpacket
	);

	Core3_id_router_003 id_router_004 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_004_src_valid),                                                                  //          .valid
		.src_data           (id_router_004_src_data),                                                                   //          .data
		.src_channel        (id_router_004_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                             //          .endofpacket
	);

	Core3_id_router_005 id_router_005 (
		.sink_ready         (mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mutex_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                               //       src.ready
		.src_valid          (id_router_005_src_valid),                                               //          .valid
		.src_data           (id_router_005_src_data),                                                //          .data
		.src_channel        (id_router_005_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                          //          .endofpacket
	);

	Core3_id_router_005 id_router_006 (
		.sink_ready         (mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mutex_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                               //       src.ready
		.src_valid          (id_router_006_src_valid),                                               //          .valid
		.src_data           (id_router_006_src_data),                                                //          .data
		.src_channel        (id_router_006_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                          //          .endofpacket
	);

	Core3_id_router_005 id_router_007 (
		.sink_ready         (mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mutex_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                               //       src.ready
		.src_valid          (id_router_007_src_valid),                                               //          .valid
		.src_data           (id_router_007_src_data),                                                //          .data
		.src_channel        (id_router_007_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                          //          .endofpacket
	);

	Core3_id_router_005 id_router_008 (
		.sink_ready         (mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mutex_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                               //       src.ready
		.src_valid          (id_router_008_src_valid),                                               //          .valid
		.src_data           (id_router_008_src_data),                                                //          .data
		.src_channel        (id_router_008_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                          //          .endofpacket
	);

	Core3_id_router_005 id_router_009 (
		.sink_ready         (mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mutex_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                               //       src.ready
		.src_valid          (id_router_009_src_valid),                                               //          .valid
		.src_data           (id_router_009_src_data),                                                //          .data
		.src_channel        (id_router_009_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                          //          .endofpacket
	);

	Core3_id_router_005 id_router_010 (
		.sink_ready         (mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mutex_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                               //       src.ready
		.src_valid          (id_router_010_src_valid),                                               //          .valid
		.src_data           (id_router_010_src_data),                                                //          .data
		.src_channel        (id_router_010_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                          //          .endofpacket
	);

	Core3_id_router_003 id_router_011 (
		.sink_ready         (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_to_1_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                   //       src.ready
		.src_valid          (id_router_011_src_valid),                                                   //          .valid
		.src_data           (id_router_011_src_data),                                                    //          .data
		.src_channel        (id_router_011_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                              //          .endofpacket
	);

	Core3_id_router_003 id_router_012 (
		.sink_ready         (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                       //       src.ready
		.src_valid          (id_router_012_src_valid),                                                       //          .valid
		.src_data           (id_router_012_src_data),                                                        //          .data
		.src_channel        (id_router_012_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                  //          .endofpacket
	);

	Core3_id_router_003 id_router_013 (
		.sink_ready         (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                   //       src.ready
		.src_valid          (id_router_013_src_valid),                                                   //          .valid
		.src_data           (id_router_013_src_data),                                                    //          .data
		.src_channel        (id_router_013_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                              //          .endofpacket
	);

	Core3_id_router_003 id_router_014 (
		.sink_ready         (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                       //       src.ready
		.src_valid          (id_router_014_src_valid),                                                       //          .valid
		.src_data           (id_router_014_src_data),                                                        //          .data
		.src_channel        (id_router_014_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                  //          .endofpacket
	);

	Core3_id_router_003 id_router_015 (
		.sink_ready         (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_1_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                        //       src.ready
		.src_valid          (id_router_015_src_valid),                                                        //          .valid
		.src_data           (id_router_015_src_data),                                                         //          .data
		.src_channel        (id_router_015_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                   //          .endofpacket
	);

	Core3_id_router_003 id_router_016 (
		.sink_ready         (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_1_to_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                    //       src.ready
		.src_valid          (id_router_016_src_valid),                                                    //          .valid
		.src_data           (id_router_016_src_data),                                                     //          .data
		.src_channel        (id_router_016_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                               //          .endofpacket
	);

	Core3_id_router_003 id_router_017 (
		.sink_ready         (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_2_to_0_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                    //       src.ready
		.src_valid          (id_router_017_src_valid),                                                    //          .valid
		.src_data           (id_router_017_src_data),                                                     //          .data
		.src_channel        (id_router_017_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                               //          .endofpacket
	);

	Core3_id_router_003 id_router_018 (
		.sink_ready         (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_2_to_0_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                        //       src.ready
		.src_valid          (id_router_018_src_valid),                                                        //          .valid
		.src_data           (id_router_018_src_data),                                                         //          .data
		.src_channel        (id_router_018_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                                   //          .endofpacket
	);

	Core3_id_router_005 id_router_019 (
		.sink_ready         (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (red_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                //       src.ready
		.src_valid          (id_router_019_src_valid),                                                //          .valid
		.src_data           (id_router_019_src_data),                                                 //          .data
		.src_channel        (id_router_019_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                           //          .endofpacket
	);

	Core3_id_router_005 id_router_020 (
		.sink_ready         (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                                  //       src.ready
		.src_valid          (id_router_020_src_valid),                                                  //          .valid
		.src_data           (id_router_020_src_data),                                                   //          .data
		.src_channel        (id_router_020_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                             //          .endofpacket
	);

	Core3_id_router_005 id_router_021 (
		.sink_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switches_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                                //       src.ready
		.src_valid          (id_router_021_src_valid),                                                //          .valid
		.src_data           (id_router_021_src_data),                                                 //          .data
		.src_channel        (id_router_021_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                           //          .endofpacket
	);

	Core3_id_router_005 id_router_022 (
		.sink_ready         (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_shared_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                                      //       src.ready
		.src_valid          (id_router_022_src_valid),                                                      //          .valid
		.src_data           (id_router_022_src_data),                                                       //          .data
		.src_channel        (id_router_022_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                                 //          .endofpacket
	);

	Core3_id_router_003 id_router_023 (
		.sink_ready         (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                                                                        //       src.ready
		.src_valid          (id_router_023_src_valid),                                                                        //          .valid
		.src_data           (id_router_023_src_data),                                                                         //          .data
		.src_channel        (id_router_023_src_channel),                                                                      //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),                                                                //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)                                                                   //          .endofpacket
	);

	Core3_id_router_003 id_router_024 (
		.sink_ready         (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                                                 //       src.ready
		.src_valid          (id_router_024_src_valid),                                                 //          .valid
		.src_data           (id_router_024_src_data),                                                  //          .data
		.src_channel        (id_router_024_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)                                            //          .endofpacket
	);

	Core3_id_router_005 id_router_025 (
		.sink_ready         (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_shared_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_025_src_ready),                                                      //       src.ready
		.src_valid          (id_router_025_src_valid),                                                      //          .valid
		.src_data           (id_router_025_src_data),                                                       //          .data
		.src_channel        (id_router_025_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_025_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_025_src_endofpacket)                                                 //          .endofpacket
	);

	Core3_id_router_026 id_router_026 (
		.sink_ready         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_1_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_026_src_ready),                                                            //       src.ready
		.src_valid          (id_router_026_src_valid),                                                            //          .valid
		.src_data           (id_router_026_src_data),                                                             //          .data
		.src_channel        (id_router_026_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_026_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_026_src_endofpacket)                                                       //          .endofpacket
	);

	Core3_id_router_026 id_router_027 (
		.sink_ready         (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_027_src_ready),                                                       //       src.ready
		.src_valid          (id_router_027_src_valid),                                                       //          .valid
		.src_data           (id_router_027_src_data),                                                        //          .data
		.src_channel        (id_router_027_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_027_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_027_src_endofpacket)                                                  //          .endofpacket
	);

	Core3_id_router_028 id_router_028 (
		.sink_ready         (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_1_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_028_src_ready),                                                 //       src.ready
		.src_valid          (id_router_028_src_valid),                                                 //          .valid
		.src_data           (id_router_028_src_data),                                                  //          .data
		.src_channel        (id_router_028_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_028_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_028_src_endofpacket)                                            //          .endofpacket
	);

	Core3_id_router_028 id_router_029 (
		.sink_ready         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_1_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_029_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_029_src_valid),                                                                  //          .valid
		.src_data           (id_router_029_src_data),                                                                   //          .data
		.src_channel        (id_router_029_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_029_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_029_src_endofpacket)                                                             //          .endofpacket
	);

	Core3_id_router_028 id_router_030 (
		.sink_ready         (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_to_1_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_030_src_ready),                                                    //       src.ready
		.src_valid          (id_router_030_src_valid),                                                    //          .valid
		.src_data           (id_router_030_src_data),                                                     //          .data
		.src_channel        (id_router_030_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_030_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_030_src_endofpacket)                                               //          .endofpacket
	);

	Core3_id_router_028 id_router_031 (
		.sink_ready         (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_031_src_ready),                                                        //       src.ready
		.src_valid          (id_router_031_src_valid),                                                        //          .valid
		.src_data           (id_router_031_src_data),                                                         //          .data
		.src_channel        (id_router_031_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_031_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_031_src_endofpacket)                                                   //          .endofpacket
	);

	Core3_id_router_028 id_router_032 (
		.sink_ready         (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_1_to_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_032_src_ready),                                                   //       src.ready
		.src_valid          (id_router_032_src_valid),                                                   //          .valid
		.src_data           (id_router_032_src_data),                                                    //          .data
		.src_channel        (id_router_032_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_032_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_032_src_endofpacket)                                              //          .endofpacket
	);

	Core3_id_router_028 id_router_033 (
		.sink_ready         (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_1_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_033_src_ready),                                                       //       src.ready
		.src_valid          (id_router_033_src_valid),                                                       //          .valid
		.src_data           (id_router_033_src_data),                                                        //          .data
		.src_channel        (id_router_033_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_033_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_033_src_endofpacket)                                                  //          .endofpacket
	);

	Core3_id_router_028 id_router_034 (
		.sink_ready         (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_1_to_2_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_034_src_ready),                                                   //       src.ready
		.src_valid          (id_router_034_src_valid),                                                   //          .valid
		.src_data           (id_router_034_src_data),                                                    //          .data
		.src_channel        (id_router_034_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_034_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_034_src_endofpacket)                                              //          .endofpacket
	);

	Core3_id_router_028 id_router_035 (
		.sink_ready         (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_1_to_2_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_035_src_ready),                                                       //       src.ready
		.src_valid          (id_router_035_src_valid),                                                       //          .valid
		.src_data           (id_router_035_src_data),                                                        //          .data
		.src_channel        (id_router_035_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_035_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_035_src_endofpacket)                                                  //          .endofpacket
	);

	Core3_id_router_028 id_router_036 (
		.sink_ready         (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_2_to_1_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_036_src_ready),                                                    //       src.ready
		.src_valid          (id_router_036_src_valid),                                                    //          .valid
		.src_data           (id_router_036_src_data),                                                     //          .data
		.src_channel        (id_router_036_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_036_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_036_src_endofpacket)                                               //          .endofpacket
	);

	Core3_id_router_028 id_router_037 (
		.sink_ready         (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_2_to_1_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_037_src_ready),                                                        //       src.ready
		.src_valid          (id_router_037_src_valid),                                                        //          .valid
		.src_data           (id_router_037_src_data),                                                         //          .data
		.src_channel        (id_router_037_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_037_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_037_src_endofpacket)                                                   //          .endofpacket
	);

	Core3_id_router_028 id_router_038 (
		.sink_ready         (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (performance_counter_1_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                             // clk_reset.reset
		.src_ready          (id_router_038_src_ready),                                                                        //       src.ready
		.src_valid          (id_router_038_src_valid),                                                                        //          .valid
		.src_data           (id_router_038_src_data),                                                                         //          .data
		.src_channel        (id_router_038_src_channel),                                                                      //          .channel
		.src_startofpacket  (id_router_038_src_startofpacket),                                                                //          .startofpacket
		.src_endofpacket    (id_router_038_src_endofpacket)                                                                   //          .endofpacket
	);

	Core3_id_router_028 id_router_039 (
		.sink_ready         (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_1_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_039_src_ready),                                                 //       src.ready
		.src_valid          (id_router_039_src_valid),                                                 //          .valid
		.src_data           (id_router_039_src_data),                                                  //          .data
		.src_channel        (id_router_039_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_039_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_039_src_endofpacket)                                            //          .endofpacket
	);

	Core3_id_router_040 id_router_040 (
		.sink_ready         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_040_src_ready),                                                            //       src.ready
		.src_valid          (id_router_040_src_valid),                                                            //          .valid
		.src_data           (id_router_040_src_data),                                                             //          .data
		.src_channel        (id_router_040_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_040_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_040_src_endofpacket)                                                       //          .endofpacket
	);

	Core3_id_router_040 id_router_041 (
		.sink_ready         (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_041_src_ready),                                                       //       src.ready
		.src_valid          (id_router_041_src_valid),                                                       //          .valid
		.src_data           (id_router_041_src_data),                                                        //          .data
		.src_channel        (id_router_041_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_041_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_041_src_endofpacket)                                                  //          .endofpacket
	);

	Core3_id_router_042 id_router_042 (
		.sink_ready         (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_042_src_ready),                                                 //       src.ready
		.src_valid          (id_router_042_src_valid),                                                 //          .valid
		.src_data           (id_router_042_src_data),                                                  //          .data
		.src_channel        (id_router_042_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_042_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_042_src_endofpacket)                                            //          .endofpacket
	);

	Core3_id_router_042 id_router_043 (
		.sink_ready         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_2_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_043_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_043_src_valid),                                                                  //          .valid
		.src_data           (id_router_043_src_data),                                                                   //          .data
		.src_channel        (id_router_043_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_043_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_043_src_endofpacket)                                                             //          .endofpacket
	);

	Core3_id_router_042 id_router_044 (
		.sink_ready         (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_044_src_ready),                                                    //       src.ready
		.src_valid          (id_router_044_src_valid),                                                    //          .valid
		.src_data           (id_router_044_src_data),                                                     //          .data
		.src_channel        (id_router_044_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_044_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_044_src_endofpacket)                                               //          .endofpacket
	);

	Core3_id_router_042 id_router_045 (
		.sink_ready         (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_045_src_ready),                                                        //       src.ready
		.src_valid          (id_router_045_src_valid),                                                        //          .valid
		.src_data           (id_router_045_src_data),                                                         //          .data
		.src_channel        (id_router_045_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_045_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_045_src_endofpacket)                                                   //          .endofpacket
	);

	Core3_id_router_042 id_router_046 (
		.sink_ready         (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_1_to_2_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_046_src_ready),                                                    //       src.ready
		.src_valid          (id_router_046_src_valid),                                                    //          .valid
		.src_data           (id_router_046_src_data),                                                     //          .data
		.src_channel        (id_router_046_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_046_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_046_src_endofpacket)                                               //          .endofpacket
	);

	Core3_id_router_042 id_router_047 (
		.sink_ready         (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_1_to_2_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_047_src_ready),                                                        //       src.ready
		.src_valid          (id_router_047_src_valid),                                                        //          .valid
		.src_data           (id_router_047_src_data),                                                         //          .data
		.src_channel        (id_router_047_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_047_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_047_src_endofpacket)                                                   //          .endofpacket
	);

	Core3_id_router_042 id_router_048 (
		.sink_ready         (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_2_to_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_048_src_ready),                                                   //       src.ready
		.src_valid          (id_router_048_src_valid),                                                   //          .valid
		.src_data           (id_router_048_src_data),                                                    //          .data
		.src_channel        (id_router_048_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_048_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_048_src_endofpacket)                                              //          .endofpacket
	);

	Core3_id_router_042 id_router_049 (
		.sink_ready         (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_2_to_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_049_src_ready),                                                       //       src.ready
		.src_valid          (id_router_049_src_valid),                                                       //          .valid
		.src_data           (id_router_049_src_data),                                                        //          .data
		.src_channel        (id_router_049_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_049_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_049_src_endofpacket)                                                  //          .endofpacket
	);

	Core3_id_router_042 id_router_050 (
		.sink_ready         (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_2_to_1_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_050_src_ready),                                                   //       src.ready
		.src_valid          (id_router_050_src_valid),                                                   //          .valid
		.src_data           (id_router_050_src_data),                                                    //          .data
		.src_channel        (id_router_050_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_050_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_050_src_endofpacket)                                              //          .endofpacket
	);

	Core3_id_router_042 id_router_051 (
		.sink_ready         (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_2_to_1_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_051_src_ready),                                                       //       src.ready
		.src_valid          (id_router_051_src_valid),                                                       //          .valid
		.src_data           (id_router_051_src_data),                                                        //          .data
		.src_channel        (id_router_051_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_051_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_051_src_endofpacket)                                                  //          .endofpacket
	);

	Core3_id_router_042 id_router_052 (
		.sink_ready         (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (performance_counter_2_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                        //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                             // clk_reset.reset
		.src_ready          (id_router_052_src_ready),                                                                        //       src.ready
		.src_valid          (id_router_052_src_valid),                                                                        //          .valid
		.src_data           (id_router_052_src_data),                                                                         //          .data
		.src_channel        (id_router_052_src_channel),                                                                      //          .channel
		.src_startofpacket  (id_router_052_src_startofpacket),                                                                //          .startofpacket
		.src_endofpacket    (id_router_052_src_endofpacket)                                                                   //          .endofpacket
	);

	Core3_id_router_042 id_router_053 (
		.sink_ready         (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_2_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_053_src_ready),                                                 //       src.ready
		.src_valid          (id_router_053_src_valid),                                                 //          .valid
		.src_data           (id_router_053_src_data),                                                  //          .data
		.src_channel        (id_router_053_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_053_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_053_src_endofpacket)                                            //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller (
		.reset_in0  (cpu_0_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                      // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller_001 (
		.reset_in0  (cpu_1_jtag_debug_module_reset_reset),    // reset_in0.reset
		.reset_in1  (~reset_reset_n),                         // reset_in1.reset
		.clk        (clk_clk),                                //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req  (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_in2  (1'b0),                                   // (terminated)
		.reset_in3  (1'b0),                                   // (terminated)
		.reset_in4  (1'b0),                                   // (terminated)
		.reset_in5  (1'b0),                                   // (terminated)
		.reset_in6  (1'b0),                                   // (terminated)
		.reset_in7  (1'b0),                                   // (terminated)
		.reset_in8  (1'b0),                                   // (terminated)
		.reset_in9  (1'b0),                                   // (terminated)
		.reset_in10 (1'b0),                                   // (terminated)
		.reset_in11 (1'b0),                                   // (terminated)
		.reset_in12 (1'b0),                                   // (terminated)
		.reset_in13 (1'b0),                                   // (terminated)
		.reset_in14 (1'b0),                                   // (terminated)
		.reset_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (4),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller_002 (
		.reset_in0  (cpu_0_jtag_debug_module_reset_reset),    // reset_in0.reset
		.reset_in1  (cpu_1_jtag_debug_module_reset_reset),    // reset_in1.reset
		.reset_in2  (cpu_2_jtag_debug_module_reset_reset),    // reset_in2.reset
		.reset_in3  (~reset_reset_n),                         // reset_in3.reset
		.clk        (clk_clk),                                //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req  (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_in4  (1'b0),                                   // (terminated)
		.reset_in5  (1'b0),                                   // (terminated)
		.reset_in6  (1'b0),                                   // (terminated)
		.reset_in7  (1'b0),                                   // (terminated)
		.reset_in8  (1'b0),                                   // (terminated)
		.reset_in9  (1'b0),                                   // (terminated)
		.reset_in10 (1'b0),                                   // (terminated)
		.reset_in11 (1'b0),                                   // (terminated)
		.reset_in12 (1'b0),                                   // (terminated)
		.reset_in13 (1'b0),                                   // (terminated)
		.reset_in14 (1'b0),                                   // (terminated)
		.reset_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller_003 (
		.reset_in0  (cpu_2_jtag_debug_module_reset_reset),    // reset_in0.reset
		.reset_in1  (~reset_reset_n),                         // reset_in1.reset
		.clk        (clk_clk),                                //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req  (rst_controller_003_reset_out_reset_req), //          .reset_req
		.reset_in2  (1'b0),                                   // (terminated)
		.reset_in3  (1'b0),                                   // (terminated)
		.reset_in4  (1'b0),                                   // (terminated)
		.reset_in5  (1'b0),                                   // (terminated)
		.reset_in6  (1'b0),                                   // (terminated)
		.reset_in7  (1'b0),                                   // (terminated)
		.reset_in8  (1'b0),                                   // (terminated)
		.reset_in9  (1'b0),                                   // (terminated)
		.reset_in10 (1'b0),                                   // (terminated)
		.reset_in11 (1'b0),                                   // (terminated)
		.reset_in12 (1'b0),                                   // (terminated)
		.reset_in13 (1'b0),                                   // (terminated)
		.reset_in14 (1'b0),                                   // (terminated)
		.reset_in15 (1'b0)                                    // (terminated)
	);

	Core3_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_001_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_001_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_001_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_001_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_001_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_001_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_001_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_001_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_001_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_001_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_001_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_001_src20_endofpacket),   //          .endofpacket
		.src21_ready         (cmd_xbar_demux_001_src21_ready),         //     src21.ready
		.src21_valid         (cmd_xbar_demux_001_src21_valid),         //          .valid
		.src21_data          (cmd_xbar_demux_001_src21_data),          //          .data
		.src21_channel       (cmd_xbar_demux_001_src21_channel),       //          .channel
		.src21_startofpacket (cmd_xbar_demux_001_src21_startofpacket), //          .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_001_src21_endofpacket),   //          .endofpacket
		.src22_ready         (cmd_xbar_demux_001_src22_ready),         //     src22.ready
		.src22_valid         (cmd_xbar_demux_001_src22_valid),         //          .valid
		.src22_data          (cmd_xbar_demux_001_src22_data),          //          .data
		.src22_channel       (cmd_xbar_demux_001_src22_channel),       //          .channel
		.src22_startofpacket (cmd_xbar_demux_001_src22_startofpacket), //          .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_001_src22_endofpacket),   //          .endofpacket
		.src23_ready         (cmd_xbar_demux_001_src23_ready),         //     src23.ready
		.src23_valid         (cmd_xbar_demux_001_src23_valid),         //          .valid
		.src23_data          (cmd_xbar_demux_001_src23_data),          //          .data
		.src23_channel       (cmd_xbar_demux_001_src23_channel),       //          .channel
		.src23_startofpacket (cmd_xbar_demux_001_src23_startofpacket), //          .startofpacket
		.src23_endofpacket   (cmd_xbar_demux_001_src23_endofpacket),   //          .endofpacket
		.src24_ready         (cmd_xbar_demux_001_src24_ready),         //     src24.ready
		.src24_valid         (cmd_xbar_demux_001_src24_valid),         //          .valid
		.src24_data          (cmd_xbar_demux_001_src24_data),          //          .data
		.src24_channel       (cmd_xbar_demux_001_src24_channel),       //          .channel
		.src24_startofpacket (cmd_xbar_demux_001_src24_startofpacket), //          .startofpacket
		.src24_endofpacket   (cmd_xbar_demux_001_src24_endofpacket),   //          .endofpacket
		.src25_ready         (cmd_xbar_demux_001_src25_ready),         //     src25.ready
		.src25_valid         (cmd_xbar_demux_001_src25_valid),         //          .valid
		.src25_data          (cmd_xbar_demux_001_src25_data),          //          .data
		.src25_channel       (cmd_xbar_demux_001_src25_channel),       //          .channel
		.src25_startofpacket (cmd_xbar_demux_001_src25_startofpacket), //          .startofpacket
		.src25_endofpacket   (cmd_xbar_demux_001_src25_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux_001 cmd_xbar_demux_002 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.sink_ready          (addr_router_002_src_ready),              //      sink.ready
		.sink_channel        (addr_router_002_src_channel),            //          .channel
		.sink_data           (addr_router_002_src_data),               //          .data
		.sink_startofpacket  (addr_router_002_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_002_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_002_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_002_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_002_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_002_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_002_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_002_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_002_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_002_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_002_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_002_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_002_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_002_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_002_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_002_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_002_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_002_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_002_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_002_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_002_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_002_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_002_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_002_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_002_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_002_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_002_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_002_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_002_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_002_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_002_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_002_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_002_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_002_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_002_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_002_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_002_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_002_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_002_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_002_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_002_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_002_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_002_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_002_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_002_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_002_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_002_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_002_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_002_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_002_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_002_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_002_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_002_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_002_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_002_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_002_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_002_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_002_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_002_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_002_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_002_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_002_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_002_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_002_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_002_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_002_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_002_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_002_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_002_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_002_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_002_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_002_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_002_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_002_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_002_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_002_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_002_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_002_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_002_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_002_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_002_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_002_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_002_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_002_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_002_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_002_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_002_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_002_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_002_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_002_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_002_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_002_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_002_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_002_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_002_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_002_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_002_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_002_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_002_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_002_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_002_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_002_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_002_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_002_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_002_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_002_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_002_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_002_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_002_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_002_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_002_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_002_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_002_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_002_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_002_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_002_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_002_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_002_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_002_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_002_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_002_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_002_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_002_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_002_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_002_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_002_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_002_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_002_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_002_src20_endofpacket),   //          .endofpacket
		.src21_ready         (cmd_xbar_demux_002_src21_ready),         //     src21.ready
		.src21_valid         (cmd_xbar_demux_002_src21_valid),         //          .valid
		.src21_data          (cmd_xbar_demux_002_src21_data),          //          .data
		.src21_channel       (cmd_xbar_demux_002_src21_channel),       //          .channel
		.src21_startofpacket (cmd_xbar_demux_002_src21_startofpacket), //          .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_002_src21_endofpacket),   //          .endofpacket
		.src22_ready         (cmd_xbar_demux_002_src22_ready),         //     src22.ready
		.src22_valid         (cmd_xbar_demux_002_src22_valid),         //          .valid
		.src22_data          (cmd_xbar_demux_002_src22_data),          //          .data
		.src22_channel       (cmd_xbar_demux_002_src22_channel),       //          .channel
		.src22_startofpacket (cmd_xbar_demux_002_src22_startofpacket), //          .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_002_src22_endofpacket),   //          .endofpacket
		.src23_ready         (cmd_xbar_demux_002_src23_ready),         //     src23.ready
		.src23_valid         (cmd_xbar_demux_002_src23_valid),         //          .valid
		.src23_data          (cmd_xbar_demux_002_src23_data),          //          .data
		.src23_channel       (cmd_xbar_demux_002_src23_channel),       //          .channel
		.src23_startofpacket (cmd_xbar_demux_002_src23_startofpacket), //          .startofpacket
		.src23_endofpacket   (cmd_xbar_demux_002_src23_endofpacket),   //          .endofpacket
		.src24_ready         (cmd_xbar_demux_002_src24_ready),         //     src24.ready
		.src24_valid         (cmd_xbar_demux_002_src24_valid),         //          .valid
		.src24_data          (cmd_xbar_demux_002_src24_data),          //          .data
		.src24_channel       (cmd_xbar_demux_002_src24_channel),       //          .channel
		.src24_startofpacket (cmd_xbar_demux_002_src24_startofpacket), //          .startofpacket
		.src24_endofpacket   (cmd_xbar_demux_002_src24_endofpacket),   //          .endofpacket
		.src25_ready         (cmd_xbar_demux_002_src25_ready),         //     src25.ready
		.src25_valid         (cmd_xbar_demux_002_src25_valid),         //          .valid
		.src25_data          (cmd_xbar_demux_002_src25_data),          //          .data
		.src25_channel       (cmd_xbar_demux_002_src25_channel),       //          .channel
		.src25_startofpacket (cmd_xbar_demux_002_src25_startofpacket), //          .startofpacket
		.src25_endofpacket   (cmd_xbar_demux_002_src25_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux cmd_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_003_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_003_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_003_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_003_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_003_src2_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux_001 cmd_xbar_demux_004 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),     // clk_reset.reset
		.sink_ready          (addr_router_004_src_ready),              //      sink.ready
		.sink_channel        (addr_router_004_src_channel),            //          .channel
		.sink_data           (addr_router_004_src_data),               //          .data
		.sink_startofpacket  (addr_router_004_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_004_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_004_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_004_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_004_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_004_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_004_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_004_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_004_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_004_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_004_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_004_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_004_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_004_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_004_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_004_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_004_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_004_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_004_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_004_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_004_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_004_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_004_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_004_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_004_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_004_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_004_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_004_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_004_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_004_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_004_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_004_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_004_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_004_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_004_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_004_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_004_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_004_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_004_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_004_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_004_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_004_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_004_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_004_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_004_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_004_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_004_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_004_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_004_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_004_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_004_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_004_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_004_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_004_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_004_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_004_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_004_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_004_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_004_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_004_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_004_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_004_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_004_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_004_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_004_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_004_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_004_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_004_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_004_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_004_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_004_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_004_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_004_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_004_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_004_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_004_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_004_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_004_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_004_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_004_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_004_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_004_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_004_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_004_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_004_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_004_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_004_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_004_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_004_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_004_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_004_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_004_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_004_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_004_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_004_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_004_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_004_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_004_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_004_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_004_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_004_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_004_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_004_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_004_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_004_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_004_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_004_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_004_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_004_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_004_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_004_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_004_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_004_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_004_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_004_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_004_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_004_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_004_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_004_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_004_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_004_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_004_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_004_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_004_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_004_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_004_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_004_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_004_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_004_src20_endofpacket),   //          .endofpacket
		.src21_ready         (cmd_xbar_demux_004_src21_ready),         //     src21.ready
		.src21_valid         (cmd_xbar_demux_004_src21_valid),         //          .valid
		.src21_data          (cmd_xbar_demux_004_src21_data),          //          .data
		.src21_channel       (cmd_xbar_demux_004_src21_channel),       //          .channel
		.src21_startofpacket (cmd_xbar_demux_004_src21_startofpacket), //          .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_004_src21_endofpacket),   //          .endofpacket
		.src22_ready         (cmd_xbar_demux_004_src22_ready),         //     src22.ready
		.src22_valid         (cmd_xbar_demux_004_src22_valid),         //          .valid
		.src22_data          (cmd_xbar_demux_004_src22_data),          //          .data
		.src22_channel       (cmd_xbar_demux_004_src22_channel),       //          .channel
		.src22_startofpacket (cmd_xbar_demux_004_src22_startofpacket), //          .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_004_src22_endofpacket),   //          .endofpacket
		.src23_ready         (cmd_xbar_demux_004_src23_ready),         //     src23.ready
		.src23_valid         (cmd_xbar_demux_004_src23_valid),         //          .valid
		.src23_data          (cmd_xbar_demux_004_src23_data),          //          .data
		.src23_channel       (cmd_xbar_demux_004_src23_channel),       //          .channel
		.src23_startofpacket (cmd_xbar_demux_004_src23_startofpacket), //          .startofpacket
		.src23_endofpacket   (cmd_xbar_demux_004_src23_endofpacket),   //          .endofpacket
		.src24_ready         (cmd_xbar_demux_004_src24_ready),         //     src24.ready
		.src24_valid         (cmd_xbar_demux_004_src24_valid),         //          .valid
		.src24_data          (cmd_xbar_demux_004_src24_data),          //          .data
		.src24_channel       (cmd_xbar_demux_004_src24_channel),       //          .channel
		.src24_startofpacket (cmd_xbar_demux_004_src24_startofpacket), //          .startofpacket
		.src24_endofpacket   (cmd_xbar_demux_004_src24_endofpacket),   //          .endofpacket
		.src25_ready         (cmd_xbar_demux_004_src25_ready),         //     src25.ready
		.src25_valid         (cmd_xbar_demux_004_src25_valid),         //          .valid
		.src25_data          (cmd_xbar_demux_004_src25_data),          //          .data
		.src25_channel       (cmd_xbar_demux_004_src25_channel),       //          .channel
		.src25_startofpacket (cmd_xbar_demux_004_src25_startofpacket), //          .startofpacket
		.src25_endofpacket   (cmd_xbar_demux_004_src25_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux cmd_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_005_src_ready),             //      sink.ready
		.sink_channel       (addr_router_005_src_channel),           //          .channel
		.sink_data          (addr_router_005_src_data),              //          .data
		.sink_startofpacket (addr_router_005_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_005_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_005_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_005_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_005_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_005_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_005_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_005_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_005_src2_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_mux_002 cmd_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (cmd_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (cmd_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_mux_005 cmd_xbar_mux_005 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src5_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src1_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src1_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src1_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_004_src1_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_mux_005 cmd_xbar_mux_006 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_006_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_006_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_006_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_006_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_006_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_006_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src6_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src6_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src6_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src6_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src2_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src2_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src2_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_004_src2_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src2_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src2_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_mux_005 cmd_xbar_mux_007 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_007_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_007_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_007_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_007_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_007_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_007_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src7_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src7_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src7_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src7_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src7_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src3_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src3_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src3_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src3_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_004_src3_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src3_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src3_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_mux_005 cmd_xbar_mux_008 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_008_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_008_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_008_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src8_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src8_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src8_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src8_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src8_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src8_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src4_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src4_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src4_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src4_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_004_src4_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src4_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src4_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_mux_005 cmd_xbar_mux_009 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_009_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_009_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_009_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_009_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_009_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_009_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src9_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src9_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src9_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src9_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src9_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src9_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src5_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src5_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src5_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src5_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src5_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src5_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src5_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src5_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src5_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_004_src5_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src5_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src5_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_mux_005 cmd_xbar_mux_010 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_010_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_010_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_010_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_010_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_010_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_010_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src10_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src6_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src6_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src6_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_002_src6_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src6_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src6_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src6_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src6_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src6_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_004_src6_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src6_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src6_endofpacket)     //          .endofpacket
	);

	Core3_cmd_xbar_mux_005 cmd_xbar_mux_019 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_019_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_019_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_019_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_019_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_019_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_019_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src19_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src19_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src19_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src19_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src19_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src19_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src7_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src7_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src7_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_002_src7_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src7_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src7_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src7_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src7_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src7_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_004_src7_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src7_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src7_endofpacket)     //          .endofpacket
	);

	Core3_cmd_xbar_mux_005 cmd_xbar_mux_020 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_020_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_020_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_020_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_020_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_020_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_020_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src20_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src20_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src20_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src20_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src20_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src20_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src8_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src8_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src8_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_002_src8_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src8_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src8_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src8_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src8_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src8_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_004_src8_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src8_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src8_endofpacket)     //          .endofpacket
	);

	Core3_cmd_xbar_mux_005 cmd_xbar_mux_021 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_021_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_021_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_021_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_021_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_021_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_021_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src21_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src21_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src21_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src21_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src21_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src21_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src9_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src9_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src9_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_002_src9_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src9_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src9_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src9_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src9_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src9_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_004_src9_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src9_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src9_endofpacket)     //          .endofpacket
	);

	Core3_cmd_xbar_mux_005 cmd_xbar_mux_022 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_022_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_022_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_022_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_022_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_022_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_022_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src22_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src22_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src22_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src22_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src22_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src22_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src10_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src10_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src10_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src10_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src10_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src10_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src10_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src10_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src10_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_004_src10_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src10_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src10_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_mux_005 cmd_xbar_mux_025 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_025_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_025_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_025_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_025_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_025_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_025_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src25_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src25_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src25_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src25_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src25_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src25_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src11_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src11_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src11_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src11_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src11_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src11_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src11_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src11_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src11_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_004_src11_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src11_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src11_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_mux cmd_xbar_mux_026 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_026_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_026_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_026_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_026_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_026_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_026_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src12_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src12_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src12_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src12_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src12_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src12_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src1_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src1_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src1_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_003_src1_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src1_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket)     //          .endofpacket
	);

	Core3_cmd_xbar_mux cmd_xbar_mux_027 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_027_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_027_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_027_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_027_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_027_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_027_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src13_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src13_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src13_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src13_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src13_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src13_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src2_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src2_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src2_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_003_src2_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src2_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src2_endofpacket)     //          .endofpacket
	);

	Core3_cmd_xbar_mux cmd_xbar_mux_040 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_040_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_040_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_040_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_040_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_040_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_040_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_004_src12_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_004_src12_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_004_src12_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_004_src12_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_004_src12_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_004_src12_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_005_src1_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_005_src1_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_005_src1_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_005_src1_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_005_src1_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_005_src1_endofpacket)     //          .endofpacket
	);

	Core3_cmd_xbar_mux cmd_xbar_mux_041 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_041_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_041_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_041_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_041_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_041_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_041_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_004_src13_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_004_src13_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_004_src13_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_004_src13_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_004_src13_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_004_src13_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_005_src2_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_005_src2_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_005_src2_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_005_src2_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_005_src2_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_005_src2_endofpacket)     //          .endofpacket
	);

	Core3_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_002_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_002_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_002_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_002_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_002_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_002_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_002_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_002_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_002_src3_endofpacket),   //          .endofpacket
		.src4_ready         (rsp_xbar_demux_002_src4_ready),         //      src4.ready
		.src4_valid         (rsp_xbar_demux_002_src4_valid),         //          .valid
		.src4_data          (rsp_xbar_demux_002_src4_data),          //          .data
		.src4_channel       (rsp_xbar_demux_002_src4_channel),       //          .channel
		.src4_startofpacket (rsp_xbar_demux_002_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (rsp_xbar_demux_002_src4_endofpacket),   //          .endofpacket
		.src5_ready         (rsp_xbar_demux_002_src5_ready),         //      src5.ready
		.src5_valid         (rsp_xbar_demux_002_src5_valid),         //          .valid
		.src5_data          (rsp_xbar_demux_002_src5_data),          //          .data
		.src5_channel       (rsp_xbar_demux_002_src5_channel),       //          .channel
		.src5_startofpacket (rsp_xbar_demux_002_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (rsp_xbar_demux_002_src5_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_005_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_005_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_005_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_005_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_005_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_005_src2_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_006_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_006_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_006_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_006_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_006_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_006_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_006_src2_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_007_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_007_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_007_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_007_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_007_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_007_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_007_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_007_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_007_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_007_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_007_src2_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_008_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_008_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_008_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_008_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_008_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_008_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_008_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_008_src2_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_009_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_009_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_009_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_009_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_009_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_009_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_009_src2_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_010_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_010_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_010_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_010_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_010_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_010_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_010_src2_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_012 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_013 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_014 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_015 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_016 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_017 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_018 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux rsp_xbar_demux_019 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_019_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_019_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_019_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_019_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_019_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_019_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_019_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_019_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_019_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_019_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_019_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_019_src2_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux rsp_xbar_demux_020 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_020_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_020_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_020_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_020_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_020_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_020_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_020_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_020_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_020_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_020_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_020_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_020_src2_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux rsp_xbar_demux_021 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_021_src_ready),               //      sink.ready
		.sink_channel       (id_router_021_src_channel),             //          .channel
		.sink_data          (id_router_021_src_data),                //          .data
		.sink_startofpacket (id_router_021_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_021_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_021_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_021_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_021_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_021_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_021_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_021_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_021_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_021_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_021_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_021_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_021_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_021_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_021_src2_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux rsp_xbar_demux_022 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_022_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_022_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_022_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_022_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_022_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_022_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_022_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_022_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_022_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_022_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_022_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_022_src2_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_023 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_023_src_ready),               //      sink.ready
		.sink_channel       (id_router_023_src_channel),             //          .channel
		.sink_data          (id_router_023_src_data),                //          .data
		.sink_startofpacket (id_router_023_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_023_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_023_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_024 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_024_src_ready),               //      sink.ready
		.sink_channel       (id_router_024_src_channel),             //          .channel
		.sink_data          (id_router_024_src_data),                //          .data
		.sink_startofpacket (id_router_024_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_024_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_024_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket)    //          .endofpacket
	);

	Core3_cmd_xbar_demux rsp_xbar_demux_025 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_025_src_ready),               //      sink.ready
		.sink_channel       (id_router_025_src_channel),             //          .channel
		.sink_data          (id_router_025_src_data),                //          .data
		.sink_startofpacket (id_router_025_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_025_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_025_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_025_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_025_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_025_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_025_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_025_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_025_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_025_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_025_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_025_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_025_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_025_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_025_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_025_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_025_src2_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux rsp_xbar_demux_026 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_026_src_ready),               //      sink.ready
		.sink_channel       (id_router_026_src_channel),             //          .channel
		.sink_data          (id_router_026_src_data),                //          .data
		.sink_startofpacket (id_router_026_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_026_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_026_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_026_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_026_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_026_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_026_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_026_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_026_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_026_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_026_src1_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux rsp_xbar_demux_027 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_027_src_ready),               //      sink.ready
		.sink_channel       (id_router_027_src_channel),             //          .channel
		.sink_data          (id_router_027_src_data),                //          .data
		.sink_startofpacket (id_router_027_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_027_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_027_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_027_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_027_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_027_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_027_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_027_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_027_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_027_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_027_src1_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_028 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_028_src_ready),               //      sink.ready
		.sink_channel       (id_router_028_src_channel),             //          .channel
		.sink_data          (id_router_028_src_data),                //          .data
		.sink_startofpacket (id_router_028_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_028_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_028_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_028_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_028_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_029 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_029_src_ready),               //      sink.ready
		.sink_channel       (id_router_029_src_channel),             //          .channel
		.sink_data          (id_router_029_src_data),                //          .data
		.sink_startofpacket (id_router_029_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_029_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_029_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_029_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_029_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_030 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_030_src_ready),               //      sink.ready
		.sink_channel       (id_router_030_src_channel),             //          .channel
		.sink_data          (id_router_030_src_data),                //          .data
		.sink_startofpacket (id_router_030_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_030_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_030_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_030_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_030_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_031 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_031_src_ready),               //      sink.ready
		.sink_channel       (id_router_031_src_channel),             //          .channel
		.sink_data          (id_router_031_src_data),                //          .data
		.sink_startofpacket (id_router_031_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_031_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_031_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_031_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_031_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_032 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_032_src_ready),               //      sink.ready
		.sink_channel       (id_router_032_src_channel),             //          .channel
		.sink_data          (id_router_032_src_data),                //          .data
		.sink_startofpacket (id_router_032_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_032_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_032_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_032_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_032_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_033 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_033_src_ready),               //      sink.ready
		.sink_channel       (id_router_033_src_channel),             //          .channel
		.sink_data          (id_router_033_src_data),                //          .data
		.sink_startofpacket (id_router_033_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_033_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_033_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_033_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_033_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_034 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_034_src_ready),               //      sink.ready
		.sink_channel       (id_router_034_src_channel),             //          .channel
		.sink_data          (id_router_034_src_data),                //          .data
		.sink_startofpacket (id_router_034_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_034_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_034_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_034_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_034_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_035 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_035_src_ready),               //      sink.ready
		.sink_channel       (id_router_035_src_channel),             //          .channel
		.sink_data          (id_router_035_src_data),                //          .data
		.sink_startofpacket (id_router_035_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_035_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_035_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_035_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_035_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_036 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_036_src_ready),               //      sink.ready
		.sink_channel       (id_router_036_src_channel),             //          .channel
		.sink_data          (id_router_036_src_data),                //          .data
		.sink_startofpacket (id_router_036_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_036_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_036_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_036_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_036_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_037 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_037_src_ready),               //      sink.ready
		.sink_channel       (id_router_037_src_channel),             //          .channel
		.sink_data          (id_router_037_src_data),                //          .data
		.sink_startofpacket (id_router_037_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_037_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_037_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_037_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_037_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_037_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_037_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_037_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_037_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_038 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_038_src_ready),               //      sink.ready
		.sink_channel       (id_router_038_src_channel),             //          .channel
		.sink_data          (id_router_038_src_data),                //          .data
		.sink_startofpacket (id_router_038_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_038_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_038_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_038_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_038_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_038_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_038_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_038_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_038_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_039 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_039_src_ready),               //      sink.ready
		.sink_channel       (id_router_039_src_channel),             //          .channel
		.sink_data          (id_router_039_src_data),                //          .data
		.sink_startofpacket (id_router_039_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_039_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_039_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_039_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_039_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_039_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_039_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_039_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_039_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux rsp_xbar_demux_040 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_040_src_ready),               //      sink.ready
		.sink_channel       (id_router_040_src_channel),             //          .channel
		.sink_data          (id_router_040_src_data),                //          .data
		.sink_startofpacket (id_router_040_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_040_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_040_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_040_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_040_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_040_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_040_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_040_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_040_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_040_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_040_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_040_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_040_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_040_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_040_src1_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux rsp_xbar_demux_041 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_041_src_ready),               //      sink.ready
		.sink_channel       (id_router_041_src_channel),             //          .channel
		.sink_data          (id_router_041_src_data),                //          .data
		.sink_startofpacket (id_router_041_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_041_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_041_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_041_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_041_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_041_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_041_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_041_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_041_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_041_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_041_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_041_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_041_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_041_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_041_src1_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_042 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_042_src_ready),               //      sink.ready
		.sink_channel       (id_router_042_src_channel),             //          .channel
		.sink_data          (id_router_042_src_data),                //          .data
		.sink_startofpacket (id_router_042_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_042_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_042_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_042_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_042_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_042_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_042_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_042_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_042_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_043 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_043_src_ready),               //      sink.ready
		.sink_channel       (id_router_043_src_channel),             //          .channel
		.sink_data          (id_router_043_src_data),                //          .data
		.sink_startofpacket (id_router_043_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_043_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_043_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_043_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_043_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_043_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_043_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_043_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_043_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_044 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_044_src_ready),               //      sink.ready
		.sink_channel       (id_router_044_src_channel),             //          .channel
		.sink_data          (id_router_044_src_data),                //          .data
		.sink_startofpacket (id_router_044_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_044_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_044_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_044_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_044_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_044_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_044_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_044_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_044_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_045 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_045_src_ready),               //      sink.ready
		.sink_channel       (id_router_045_src_channel),             //          .channel
		.sink_data          (id_router_045_src_data),                //          .data
		.sink_startofpacket (id_router_045_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_045_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_045_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_045_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_045_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_045_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_045_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_045_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_045_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_046 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_046_src_ready),               //      sink.ready
		.sink_channel       (id_router_046_src_channel),             //          .channel
		.sink_data          (id_router_046_src_data),                //          .data
		.sink_startofpacket (id_router_046_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_046_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_046_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_046_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_046_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_046_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_046_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_046_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_046_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_047 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_047_src_ready),               //      sink.ready
		.sink_channel       (id_router_047_src_channel),             //          .channel
		.sink_data          (id_router_047_src_data),                //          .data
		.sink_startofpacket (id_router_047_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_047_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_047_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_047_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_047_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_047_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_047_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_047_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_047_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_048 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_048_src_ready),               //      sink.ready
		.sink_channel       (id_router_048_src_channel),             //          .channel
		.sink_data          (id_router_048_src_data),                //          .data
		.sink_startofpacket (id_router_048_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_048_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_048_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_048_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_048_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_048_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_048_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_048_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_048_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_049 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_049_src_ready),               //      sink.ready
		.sink_channel       (id_router_049_src_channel),             //          .channel
		.sink_data          (id_router_049_src_data),                //          .data
		.sink_startofpacket (id_router_049_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_049_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_049_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_049_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_049_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_049_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_049_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_049_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_049_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_050 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_050_src_ready),               //      sink.ready
		.sink_channel       (id_router_050_src_channel),             //          .channel
		.sink_data          (id_router_050_src_data),                //          .data
		.sink_startofpacket (id_router_050_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_050_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_050_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_050_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_050_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_050_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_050_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_050_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_050_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_051 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_051_src_ready),               //      sink.ready
		.sink_channel       (id_router_051_src_channel),             //          .channel
		.sink_data          (id_router_051_src_data),                //          .data
		.sink_startofpacket (id_router_051_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_051_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_051_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_051_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_051_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_051_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_051_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_051_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_051_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_052 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_052_src_ready),               //      sink.ready
		.sink_channel       (id_router_052_src_channel),             //          .channel
		.sink_data          (id_router_052_src_data),                //          .data
		.sink_startofpacket (id_router_052_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_052_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_052_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_052_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_052_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_052_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_052_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_052_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_052_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_demux_003 rsp_xbar_demux_053 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_053_src_ready),               //      sink.ready
		.sink_channel       (id_router_053_src_channel),             //          .channel
		.sink_data          (id_router_053_src_data),                //          .data
		.sink_startofpacket (id_router_053_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_053_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_053_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_053_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_053_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_053_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_053_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_053_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_053_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_020_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_021_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink22_ready         (rsp_xbar_demux_022_src0_ready),         //    sink22.ready
		.sink22_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink22_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink22_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.sink22_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink22_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.sink23_ready         (rsp_xbar_demux_023_src0_ready),         //    sink23.ready
		.sink23_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink23_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink23_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.sink23_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink23_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.sink24_ready         (rsp_xbar_demux_024_src0_ready),         //    sink24.ready
		.sink24_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink24_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink24_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.sink24_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink24_endofpacket   (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.sink25_ready         (rsp_xbar_demux_025_src0_ready),         //    sink25.ready
		.sink25_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.sink25_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.sink25_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.sink25_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.sink25_endofpacket   (rsp_xbar_demux_025_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_mux_001 rsp_xbar_mux_002 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_002_src2_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_002_src2_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_002_src2_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_002_src2_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_005_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_005_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_005_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_005_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_006_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_006_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_006_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_006_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_007_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_007_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_007_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_007_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_007_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_008_src1_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_008_src1_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_008_src1_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_008_src1_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_008_src1_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_009_src1_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_009_src1_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_009_src1_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_009_src1_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_009_src1_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_010_src1_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_010_src1_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_010_src1_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_010_src1_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_019_src1_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_019_src1_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_019_src1_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_019_src1_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_019_src1_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_019_src1_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_020_src1_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_020_src1_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_020_src1_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_020_src1_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_020_src1_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_020_src1_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_021_src1_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_021_src1_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_021_src1_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_021_src1_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_021_src1_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_021_src1_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_022_src1_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_022_src1_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_022_src1_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_022_src1_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_022_src1_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_022_src1_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_025_src1_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_025_src1_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_025_src1_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_025_src1_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_025_src1_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_025_src1_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_026_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_026_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_027_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_027_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_028_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_028_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_029_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_029_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_030_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_030_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_031_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_031_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_032_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_032_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_033_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_033_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_034_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_034_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_035_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_035_src0_endofpacket),   //          .endofpacket
		.sink22_ready         (rsp_xbar_demux_036_src0_ready),         //    sink22.ready
		.sink22_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.sink22_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.sink22_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.sink22_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.sink22_endofpacket   (rsp_xbar_demux_036_src0_endofpacket),   //          .endofpacket
		.sink23_ready         (rsp_xbar_demux_037_src0_ready),         //    sink23.ready
		.sink23_valid         (rsp_xbar_demux_037_src0_valid),         //          .valid
		.sink23_channel       (rsp_xbar_demux_037_src0_channel),       //          .channel
		.sink23_data          (rsp_xbar_demux_037_src0_data),          //          .data
		.sink23_startofpacket (rsp_xbar_demux_037_src0_startofpacket), //          .startofpacket
		.sink23_endofpacket   (rsp_xbar_demux_037_src0_endofpacket),   //          .endofpacket
		.sink24_ready         (rsp_xbar_demux_038_src0_ready),         //    sink24.ready
		.sink24_valid         (rsp_xbar_demux_038_src0_valid),         //          .valid
		.sink24_channel       (rsp_xbar_demux_038_src0_channel),       //          .channel
		.sink24_data          (rsp_xbar_demux_038_src0_data),          //          .data
		.sink24_startofpacket (rsp_xbar_demux_038_src0_startofpacket), //          .startofpacket
		.sink24_endofpacket   (rsp_xbar_demux_038_src0_endofpacket),   //          .endofpacket
		.sink25_ready         (rsp_xbar_demux_039_src0_ready),         //    sink25.ready
		.sink25_valid         (rsp_xbar_demux_039_src0_valid),         //          .valid
		.sink25_channel       (rsp_xbar_demux_039_src0_channel),       //          .channel
		.sink25_data          (rsp_xbar_demux_039_src0_data),          //          .data
		.sink25_startofpacket (rsp_xbar_demux_039_src0_startofpacket), //          .startofpacket
		.sink25_endofpacket   (rsp_xbar_demux_039_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_mux rsp_xbar_mux_003 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_003_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_003_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_002_src3_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_002_src3_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_002_src3_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_002_src3_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_002_src3_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_026_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_026_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_026_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_026_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_026_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_026_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_027_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_027_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_027_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_027_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_027_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_027_src1_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_mux_001 rsp_xbar_mux_004 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_004_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_004_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_004_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_002_src4_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_002_src4_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_002_src4_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_002_src4_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_002_src4_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_002_src4_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_005_src2_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_005_src2_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_005_src2_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_005_src2_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_005_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_005_src2_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_006_src2_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_006_src2_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_006_src2_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_006_src2_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_006_src2_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_006_src2_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_007_src2_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_007_src2_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_007_src2_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_007_src2_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_007_src2_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_007_src2_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_008_src2_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_008_src2_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_008_src2_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_008_src2_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_008_src2_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_008_src2_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_009_src2_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_009_src2_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_009_src2_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_009_src2_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_009_src2_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_009_src2_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_010_src2_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_010_src2_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_010_src2_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_010_src2_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_010_src2_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_010_src2_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_019_src2_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_019_src2_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_019_src2_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_019_src2_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_019_src2_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_019_src2_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_020_src2_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_020_src2_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_020_src2_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_020_src2_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_020_src2_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_020_src2_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_021_src2_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_021_src2_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_021_src2_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_021_src2_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_021_src2_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_021_src2_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_022_src2_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_022_src2_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_022_src2_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_022_src2_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_022_src2_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_022_src2_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_025_src2_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_025_src2_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_025_src2_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_025_src2_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_025_src2_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_025_src2_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_040_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_040_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_040_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_040_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_040_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_040_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_041_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_041_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_041_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_041_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_041_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_041_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_042_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_042_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_042_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_042_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_042_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_042_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_043_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_043_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_043_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_043_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_043_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_043_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_044_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_044_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_044_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_044_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_044_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_044_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_045_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_045_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_045_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_045_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_045_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_045_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_046_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_046_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_046_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_046_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_046_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_046_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_047_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_047_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_047_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_047_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_047_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_047_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_048_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_048_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_048_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_048_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_048_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_048_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_049_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_049_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_049_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_049_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_049_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_049_src0_endofpacket),   //          .endofpacket
		.sink22_ready         (rsp_xbar_demux_050_src0_ready),         //    sink22.ready
		.sink22_valid         (rsp_xbar_demux_050_src0_valid),         //          .valid
		.sink22_channel       (rsp_xbar_demux_050_src0_channel),       //          .channel
		.sink22_data          (rsp_xbar_demux_050_src0_data),          //          .data
		.sink22_startofpacket (rsp_xbar_demux_050_src0_startofpacket), //          .startofpacket
		.sink22_endofpacket   (rsp_xbar_demux_050_src0_endofpacket),   //          .endofpacket
		.sink23_ready         (rsp_xbar_demux_051_src0_ready),         //    sink23.ready
		.sink23_valid         (rsp_xbar_demux_051_src0_valid),         //          .valid
		.sink23_channel       (rsp_xbar_demux_051_src0_channel),       //          .channel
		.sink23_data          (rsp_xbar_demux_051_src0_data),          //          .data
		.sink23_startofpacket (rsp_xbar_demux_051_src0_startofpacket), //          .startofpacket
		.sink23_endofpacket   (rsp_xbar_demux_051_src0_endofpacket),   //          .endofpacket
		.sink24_ready         (rsp_xbar_demux_052_src0_ready),         //    sink24.ready
		.sink24_valid         (rsp_xbar_demux_052_src0_valid),         //          .valid
		.sink24_channel       (rsp_xbar_demux_052_src0_channel),       //          .channel
		.sink24_data          (rsp_xbar_demux_052_src0_data),          //          .data
		.sink24_startofpacket (rsp_xbar_demux_052_src0_startofpacket), //          .startofpacket
		.sink24_endofpacket   (rsp_xbar_demux_052_src0_endofpacket),   //          .endofpacket
		.sink25_ready         (rsp_xbar_demux_053_src0_ready),         //    sink25.ready
		.sink25_valid         (rsp_xbar_demux_053_src0_valid),         //          .valid
		.sink25_channel       (rsp_xbar_demux_053_src0_channel),       //          .channel
		.sink25_data          (rsp_xbar_demux_053_src0_data),          //          .data
		.sink25_startofpacket (rsp_xbar_demux_053_src0_startofpacket), //          .startofpacket
		.sink25_endofpacket   (rsp_xbar_demux_053_src0_endofpacket)    //          .endofpacket
	);

	Core3_rsp_xbar_mux rsp_xbar_mux_005 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_005_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_005_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_002_src5_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_002_src5_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_002_src5_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_002_src5_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_002_src5_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_002_src5_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_040_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_040_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_040_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_040_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_040_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_040_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_041_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_041_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_041_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_041_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_041_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_041_src1_endofpacket)    //          .endofpacket
	);

	Core3_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (cpu_0_d_irq_irq)                 //    sender.irq
	);

	Core3_irq_mapper irq_mapper_001 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_001_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (cpu_1_d_irq_irq)                     //    sender.irq
	);

	Core3_irq_mapper irq_mapper_002 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_003_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_002_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_002_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_002_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (cpu_2_d_irq_irq)                     //    sender.irq
	);

endmodule
